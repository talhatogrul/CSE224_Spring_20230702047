magic
tech sky130A
magscale 1 2
timestamp 1745598869
<< viali >>
rect 4997 9129 5031 9163
rect 2927 9061 2961 9095
rect 5365 9061 5399 9095
rect 1409 8925 1443 8959
rect 1685 8925 1719 8959
rect 2789 8925 2823 8959
rect 3065 8925 3099 8959
rect 3249 8925 3283 8959
rect 4813 8925 4847 8959
rect 5181 8925 5215 8959
rect 1593 8789 1627 8823
rect 1869 8789 1903 8823
rect 3249 8789 3283 8823
rect 3525 8585 3559 8619
rect 2697 8449 2731 8483
rect 2973 8449 3007 8483
rect 3341 8449 3375 8483
rect 3893 8449 3927 8483
rect 5089 8449 5123 8483
rect 5273 8449 5307 8483
rect 2789 8381 2823 8415
rect 3709 8381 3743 8415
rect 4077 8381 4111 8415
rect 3157 8313 3191 8347
rect 5089 8313 5123 8347
rect 2789 8245 2823 8279
rect 2053 8041 2087 8075
rect 1777 7973 1811 8007
rect 1593 7837 1627 7871
rect 1777 7837 1811 7871
rect 1869 7837 1903 7871
rect 5181 7837 5215 7871
rect 5365 7701 5399 7735
rect 3157 7497 3191 7531
rect 3341 7361 3375 7395
rect 3433 7361 3467 7395
rect 4077 7361 4111 7395
rect 3893 7293 3927 7327
rect 4261 7157 4295 7191
rect 5089 6885 5123 6919
rect 1409 6749 1443 6783
rect 4813 6681 4847 6715
rect 1593 6613 1627 6647
rect 5273 6613 5307 6647
rect 5365 6409 5399 6443
rect 5181 6273 5215 6307
rect 2881 5797 2915 5831
rect 2421 5729 2455 5763
rect 3893 5729 3927 5763
rect 2513 5661 2547 5695
rect 3801 5661 3835 5695
rect 3985 5661 4019 5695
rect 1593 5321 1627 5355
rect 5089 5321 5123 5355
rect 1409 5185 1443 5219
rect 2789 5185 2823 5219
rect 3065 5185 3099 5219
rect 4905 5185 4939 5219
rect 5181 5185 5215 5219
rect 2973 5117 3007 5151
rect 3065 4981 3099 5015
rect 3249 4981 3283 5015
rect 5365 4981 5399 5015
rect 1409 4097 1443 4131
rect 4905 4097 4939 4131
rect 5181 4097 5215 4131
rect 1593 3961 1627 3995
rect 4721 3893 4755 3927
rect 5365 3893 5399 3927
rect 4629 3553 4663 3587
rect 5089 3553 5123 3587
rect 4721 3485 4755 3519
rect 4905 3145 4939 3179
rect 4353 3077 4387 3111
rect 4261 3009 4295 3043
rect 4445 3009 4479 3043
rect 5089 3009 5123 3043
rect 5273 3009 5307 3043
rect 5365 3009 5399 3043
rect 5181 2873 5215 2907
rect 1869 2601 1903 2635
rect 1593 2533 1627 2567
rect 4353 2533 4387 2567
rect 4077 2465 4111 2499
rect 1409 2397 1443 2431
rect 1685 2397 1719 2431
rect 3985 2397 4019 2431
rect 4629 2397 4663 2431
rect 5089 2397 5123 2431
rect 5457 2329 5491 2363
rect 4813 2261 4847 2295
<< metal1 >>
rect 1104 9274 5796 9296
rect 1104 9222 1950 9274
rect 2002 9222 2014 9274
rect 2066 9222 2078 9274
rect 2130 9222 2142 9274
rect 2194 9222 2206 9274
rect 2258 9222 5796 9274
rect 1104 9200 5796 9222
rect 4982 9120 4988 9172
rect 5040 9120 5046 9172
rect 2915 9095 2973 9101
rect 2915 9061 2927 9095
rect 2961 9092 2973 9095
rect 3050 9092 3056 9104
rect 2961 9064 3056 9092
rect 2961 9061 2973 9064
rect 2915 9055 2973 9061
rect 3050 9052 3056 9064
rect 3108 9052 3114 9104
rect 5350 9052 5356 9104
rect 5408 9052 5414 9104
rect 3418 9024 3424 9036
rect 2792 8996 3424 9024
rect 1394 8916 1400 8968
rect 1452 8916 1458 8968
rect 2792 8965 2820 8996
rect 3418 8984 3424 8996
rect 3476 8984 3482 9036
rect 1673 8959 1731 8965
rect 1673 8925 1685 8959
rect 1719 8925 1731 8959
rect 1673 8919 1731 8925
rect 2777 8959 2835 8965
rect 2777 8925 2789 8959
rect 2823 8925 2835 8959
rect 2777 8919 2835 8925
rect 3053 8959 3111 8965
rect 3053 8925 3065 8959
rect 3099 8925 3111 8959
rect 3053 8919 3111 8925
rect 842 8848 848 8900
rect 900 8888 906 8900
rect 1688 8888 1716 8919
rect 900 8860 1716 8888
rect 3068 8888 3096 8919
rect 3142 8916 3148 8968
rect 3200 8956 3206 8968
rect 3237 8959 3295 8965
rect 3237 8956 3249 8959
rect 3200 8928 3249 8956
rect 3200 8916 3206 8928
rect 3237 8925 3249 8928
rect 3283 8925 3295 8959
rect 3237 8919 3295 8925
rect 3510 8916 3516 8968
rect 3568 8956 3574 8968
rect 4801 8959 4859 8965
rect 4801 8956 4813 8959
rect 3568 8928 4813 8956
rect 3568 8916 3574 8928
rect 4801 8925 4813 8928
rect 4847 8925 4859 8959
rect 4801 8919 4859 8925
rect 5166 8916 5172 8968
rect 5224 8916 5230 8968
rect 4338 8888 4344 8900
rect 3068 8860 4344 8888
rect 900 8848 906 8860
rect 4338 8848 4344 8860
rect 4396 8848 4402 8900
rect 1578 8780 1584 8832
rect 1636 8780 1642 8832
rect 1857 8823 1915 8829
rect 1857 8789 1869 8823
rect 1903 8820 1915 8823
rect 2958 8820 2964 8832
rect 1903 8792 2964 8820
rect 1903 8789 1915 8792
rect 1857 8783 1915 8789
rect 2958 8780 2964 8792
rect 3016 8780 3022 8832
rect 3237 8823 3295 8829
rect 3237 8789 3249 8823
rect 3283 8820 3295 8823
rect 3970 8820 3976 8832
rect 3283 8792 3976 8820
rect 3283 8789 3295 8792
rect 3237 8783 3295 8789
rect 3970 8780 3976 8792
rect 4028 8780 4034 8832
rect 1104 8730 5796 8752
rect 1104 8678 2610 8730
rect 2662 8678 2674 8730
rect 2726 8678 2738 8730
rect 2790 8678 2802 8730
rect 2854 8678 2866 8730
rect 2918 8678 5796 8730
rect 1104 8656 5796 8678
rect 3510 8576 3516 8628
rect 3568 8576 3574 8628
rect 3712 8520 5304 8548
rect 2406 8440 2412 8492
rect 2464 8480 2470 8492
rect 2685 8483 2743 8489
rect 2685 8480 2697 8483
rect 2464 8452 2697 8480
rect 2464 8440 2470 8452
rect 2685 8449 2697 8452
rect 2731 8449 2743 8483
rect 2685 8443 2743 8449
rect 2958 8440 2964 8492
rect 3016 8440 3022 8492
rect 3326 8480 3332 8492
rect 3068 8452 3332 8480
rect 2774 8372 2780 8424
rect 2832 8372 2838 8424
rect 1578 8304 1584 8356
rect 1636 8344 1642 8356
rect 3068 8344 3096 8452
rect 3326 8440 3332 8452
rect 3384 8440 3390 8492
rect 3418 8372 3424 8424
rect 3476 8412 3482 8424
rect 3712 8421 3740 8520
rect 3881 8483 3939 8489
rect 3881 8449 3893 8483
rect 3927 8480 3939 8483
rect 4338 8480 4344 8492
rect 3927 8452 4344 8480
rect 3927 8449 3939 8452
rect 3881 8443 3939 8449
rect 3697 8415 3755 8421
rect 3697 8412 3709 8415
rect 3476 8384 3709 8412
rect 3476 8372 3482 8384
rect 3697 8381 3709 8384
rect 3743 8381 3755 8415
rect 3697 8375 3755 8381
rect 1636 8316 3096 8344
rect 3145 8347 3203 8353
rect 1636 8304 1642 8316
rect 2792 8285 2820 8316
rect 3145 8313 3157 8347
rect 3191 8344 3203 8347
rect 3896 8344 3924 8443
rect 4338 8440 4344 8452
rect 4396 8480 4402 8492
rect 5276 8489 5304 8520
rect 5077 8483 5135 8489
rect 5077 8480 5089 8483
rect 4396 8452 5089 8480
rect 4396 8440 4402 8452
rect 5077 8449 5089 8452
rect 5123 8449 5135 8483
rect 5077 8443 5135 8449
rect 5261 8483 5319 8489
rect 5261 8449 5273 8483
rect 5307 8449 5319 8483
rect 5261 8443 5319 8449
rect 4062 8372 4068 8424
rect 4120 8372 4126 8424
rect 3191 8316 3924 8344
rect 3191 8313 3203 8316
rect 3145 8307 3203 8313
rect 4430 8304 4436 8356
rect 4488 8344 4494 8356
rect 5077 8347 5135 8353
rect 5077 8344 5089 8347
rect 4488 8316 5089 8344
rect 4488 8304 4494 8316
rect 5077 8313 5089 8316
rect 5123 8313 5135 8347
rect 5077 8307 5135 8313
rect 2777 8279 2835 8285
rect 2777 8245 2789 8279
rect 2823 8245 2835 8279
rect 2777 8239 2835 8245
rect 1104 8186 5796 8208
rect 1104 8134 1950 8186
rect 2002 8134 2014 8186
rect 2066 8134 2078 8186
rect 2130 8134 2142 8186
rect 2194 8134 2206 8186
rect 2258 8134 5796 8186
rect 1104 8112 5796 8134
rect 2041 8075 2099 8081
rect 2041 8041 2053 8075
rect 2087 8072 2099 8075
rect 2498 8072 2504 8084
rect 2087 8044 2504 8072
rect 2087 8041 2099 8044
rect 2041 8035 2099 8041
rect 2498 8032 2504 8044
rect 2556 8072 2562 8084
rect 2774 8072 2780 8084
rect 2556 8044 2780 8072
rect 2556 8032 2562 8044
rect 2774 8032 2780 8044
rect 2832 8032 2838 8084
rect 1765 8007 1823 8013
rect 1765 7973 1777 8007
rect 1811 8004 1823 8007
rect 5166 8004 5172 8016
rect 1811 7976 5172 8004
rect 1811 7973 1823 7976
rect 1765 7967 1823 7973
rect 5166 7964 5172 7976
rect 5224 7964 5230 8016
rect 1578 7828 1584 7880
rect 1636 7828 1642 7880
rect 1762 7828 1768 7880
rect 1820 7828 1826 7880
rect 1857 7871 1915 7877
rect 1857 7837 1869 7871
rect 1903 7837 1915 7871
rect 1857 7831 1915 7837
rect 934 7760 940 7812
rect 992 7800 998 7812
rect 1872 7800 1900 7831
rect 4154 7828 4160 7880
rect 4212 7868 4218 7880
rect 5169 7871 5227 7877
rect 5169 7868 5181 7871
rect 4212 7840 5181 7868
rect 4212 7828 4218 7840
rect 5169 7837 5181 7840
rect 5215 7837 5227 7871
rect 5169 7831 5227 7837
rect 992 7772 1900 7800
rect 992 7760 998 7772
rect 5350 7692 5356 7744
rect 5408 7692 5414 7744
rect 1104 7642 5796 7664
rect 1104 7590 2610 7642
rect 2662 7590 2674 7642
rect 2726 7590 2738 7642
rect 2790 7590 2802 7642
rect 2854 7590 2866 7642
rect 2918 7590 5796 7642
rect 1104 7568 5796 7590
rect 1762 7488 1768 7540
rect 1820 7528 1826 7540
rect 3145 7531 3203 7537
rect 3145 7528 3157 7531
rect 1820 7500 3157 7528
rect 1820 7488 1826 7500
rect 3145 7497 3157 7500
rect 3191 7497 3203 7531
rect 3145 7491 3203 7497
rect 2958 7420 2964 7472
rect 3016 7460 3022 7472
rect 3878 7460 3884 7472
rect 3016 7432 3884 7460
rect 3016 7420 3022 7432
rect 3326 7352 3332 7404
rect 3384 7352 3390 7404
rect 3436 7401 3464 7432
rect 3878 7420 3884 7432
rect 3936 7420 3942 7472
rect 3421 7395 3479 7401
rect 3421 7361 3433 7395
rect 3467 7361 3479 7395
rect 3421 7355 3479 7361
rect 3970 7352 3976 7404
rect 4028 7392 4034 7404
rect 4065 7395 4123 7401
rect 4065 7392 4077 7395
rect 4028 7364 4077 7392
rect 4028 7352 4034 7364
rect 4065 7361 4077 7364
rect 4111 7361 4123 7395
rect 4065 7355 4123 7361
rect 3344 7324 3372 7352
rect 3786 7324 3792 7336
rect 3344 7296 3792 7324
rect 3786 7284 3792 7296
rect 3844 7284 3850 7336
rect 3881 7327 3939 7333
rect 3881 7293 3893 7327
rect 3927 7293 3939 7327
rect 3881 7287 3939 7293
rect 3234 7216 3240 7268
rect 3292 7256 3298 7268
rect 3896 7256 3924 7287
rect 3292 7228 3924 7256
rect 3292 7216 3298 7228
rect 4246 7148 4252 7200
rect 4304 7148 4310 7200
rect 1104 7098 5796 7120
rect 1104 7046 1950 7098
rect 2002 7046 2014 7098
rect 2066 7046 2078 7098
rect 2130 7046 2142 7098
rect 2194 7046 2206 7098
rect 2258 7046 5796 7098
rect 1104 7024 5796 7046
rect 5077 6919 5135 6925
rect 5077 6885 5089 6919
rect 5123 6914 5135 6919
rect 5123 6886 5157 6914
rect 5123 6885 5135 6886
rect 5077 6879 5135 6885
rect 4338 6808 4344 6860
rect 4396 6848 4402 6860
rect 5092 6848 5120 6879
rect 4396 6820 5120 6848
rect 4396 6808 4402 6820
rect 842 6740 848 6792
rect 900 6780 906 6792
rect 1397 6783 1455 6789
rect 1397 6780 1409 6783
rect 900 6752 1409 6780
rect 900 6740 906 6752
rect 1397 6749 1409 6752
rect 1443 6749 1455 6783
rect 5442 6780 5448 6792
rect 1397 6743 1455 6749
rect 3160 6752 5448 6780
rect 1581 6647 1639 6653
rect 1581 6613 1593 6647
rect 1627 6644 1639 6647
rect 2406 6644 2412 6656
rect 1627 6616 2412 6644
rect 1627 6613 1639 6616
rect 1581 6607 1639 6613
rect 2406 6604 2412 6616
rect 2464 6644 2470 6656
rect 3160 6644 3188 6752
rect 5442 6740 5448 6752
rect 5500 6740 5506 6792
rect 4798 6672 4804 6724
rect 4856 6672 4862 6724
rect 2464 6616 3188 6644
rect 2464 6604 2470 6616
rect 4890 6604 4896 6656
rect 4948 6644 4954 6656
rect 5261 6647 5319 6653
rect 5261 6644 5273 6647
rect 4948 6616 5273 6644
rect 4948 6604 4954 6616
rect 5261 6613 5273 6616
rect 5307 6613 5319 6647
rect 5261 6607 5319 6613
rect 1104 6554 5796 6576
rect 1104 6502 2610 6554
rect 2662 6502 2674 6554
rect 2726 6502 2738 6554
rect 2790 6502 2802 6554
rect 2854 6502 2866 6554
rect 2918 6502 5796 6554
rect 1104 6480 5796 6502
rect 5350 6400 5356 6452
rect 5408 6400 5414 6452
rect 5166 6264 5172 6316
rect 5224 6264 5230 6316
rect 1104 6010 5796 6032
rect 1104 5958 1950 6010
rect 2002 5958 2014 6010
rect 2066 5958 2078 6010
rect 2130 5958 2142 6010
rect 2194 5958 2206 6010
rect 2258 5958 5796 6010
rect 1104 5936 5796 5958
rect 2869 5831 2927 5837
rect 2869 5797 2881 5831
rect 2915 5828 2927 5831
rect 4154 5828 4160 5840
rect 2915 5800 4160 5828
rect 2915 5797 2927 5800
rect 2869 5791 2927 5797
rect 4154 5788 4160 5800
rect 4212 5788 4218 5840
rect 1578 5720 1584 5772
rect 1636 5760 1642 5772
rect 2409 5763 2467 5769
rect 2409 5760 2421 5763
rect 1636 5732 2421 5760
rect 1636 5720 1642 5732
rect 2409 5729 2421 5732
rect 2455 5760 2467 5763
rect 3881 5763 3939 5769
rect 3881 5760 3893 5763
rect 2455 5732 3893 5760
rect 2455 5729 2467 5732
rect 2409 5723 2467 5729
rect 3881 5729 3893 5732
rect 3927 5729 3939 5763
rect 3881 5723 3939 5729
rect 2498 5652 2504 5704
rect 2556 5652 2562 5704
rect 3786 5652 3792 5704
rect 3844 5652 3850 5704
rect 3970 5652 3976 5704
rect 4028 5652 4034 5704
rect 2516 5624 2544 5652
rect 5258 5624 5264 5636
rect 2516 5596 5264 5624
rect 5258 5584 5264 5596
rect 5316 5584 5322 5636
rect 1104 5466 5796 5488
rect 1104 5414 2610 5466
rect 2662 5414 2674 5466
rect 2726 5414 2738 5466
rect 2790 5414 2802 5466
rect 2854 5414 2866 5466
rect 2918 5414 5796 5466
rect 1104 5392 5796 5414
rect 1581 5355 1639 5361
rect 1581 5321 1593 5355
rect 1627 5352 1639 5355
rect 5077 5355 5135 5361
rect 1627 5324 3096 5352
rect 1627 5321 1639 5324
rect 1581 5315 1639 5321
rect 842 5176 848 5228
rect 900 5216 906 5228
rect 3068 5225 3096 5324
rect 5077 5321 5089 5355
rect 5123 5352 5135 5355
rect 5166 5352 5172 5364
rect 5123 5324 5172 5352
rect 5123 5321 5135 5324
rect 5077 5315 5135 5321
rect 5166 5312 5172 5324
rect 5224 5312 5230 5364
rect 1397 5219 1455 5225
rect 1397 5216 1409 5219
rect 900 5188 1409 5216
rect 900 5176 906 5188
rect 1397 5185 1409 5188
rect 1443 5185 1455 5219
rect 1397 5179 1455 5185
rect 2777 5219 2835 5225
rect 2777 5185 2789 5219
rect 2823 5185 2835 5219
rect 2777 5179 2835 5185
rect 3053 5219 3111 5225
rect 3053 5185 3065 5219
rect 3099 5216 3111 5219
rect 3326 5216 3332 5228
rect 3099 5188 3332 5216
rect 3099 5185 3111 5188
rect 3053 5179 3111 5185
rect 2792 5080 2820 5179
rect 3326 5176 3332 5188
rect 3384 5176 3390 5228
rect 4890 5176 4896 5228
rect 4948 5176 4954 5228
rect 4982 5176 4988 5228
rect 5040 5216 5046 5228
rect 5169 5219 5227 5225
rect 5169 5216 5181 5219
rect 5040 5188 5181 5216
rect 5040 5176 5046 5188
rect 5169 5185 5181 5188
rect 5215 5185 5227 5219
rect 5169 5179 5227 5185
rect 2958 5108 2964 5160
rect 3016 5148 3022 5160
rect 3142 5148 3148 5160
rect 3016 5120 3148 5148
rect 3016 5108 3022 5120
rect 3142 5108 3148 5120
rect 3200 5108 3206 5160
rect 4338 5080 4344 5092
rect 2792 5052 4344 5080
rect 4338 5040 4344 5052
rect 4396 5040 4402 5092
rect 3050 4972 3056 5024
rect 3108 4972 3114 5024
rect 3234 4972 3240 5024
rect 3292 4972 3298 5024
rect 5350 4972 5356 5024
rect 5408 4972 5414 5024
rect 1104 4922 5796 4944
rect 1104 4870 1950 4922
rect 2002 4870 2014 4922
rect 2066 4870 2078 4922
rect 2130 4870 2142 4922
rect 2194 4870 2206 4922
rect 2258 4870 5796 4922
rect 1104 4848 5796 4870
rect 1104 4378 5796 4400
rect 1104 4326 2610 4378
rect 2662 4326 2674 4378
rect 2726 4326 2738 4378
rect 2790 4326 2802 4378
rect 2854 4326 2866 4378
rect 2918 4326 5796 4378
rect 1104 4304 5796 4326
rect 842 4088 848 4140
rect 900 4128 906 4140
rect 1397 4131 1455 4137
rect 1397 4128 1409 4131
rect 900 4100 1409 4128
rect 900 4088 906 4100
rect 1397 4097 1409 4100
rect 1443 4097 1455 4131
rect 1397 4091 1455 4097
rect 4246 4088 4252 4140
rect 4304 4128 4310 4140
rect 4893 4131 4951 4137
rect 4893 4128 4905 4131
rect 4304 4100 4905 4128
rect 4304 4088 4310 4100
rect 4893 4097 4905 4100
rect 4939 4097 4951 4131
rect 4893 4091 4951 4097
rect 5166 4088 5172 4140
rect 5224 4088 5230 4140
rect 1581 3995 1639 4001
rect 1581 3961 1593 3995
rect 1627 3992 1639 3995
rect 3050 3992 3056 4004
rect 1627 3964 3056 3992
rect 1627 3961 1639 3964
rect 1581 3955 1639 3961
rect 3050 3952 3056 3964
rect 3108 3952 3114 4004
rect 4614 3884 4620 3936
rect 4672 3924 4678 3936
rect 4709 3927 4767 3933
rect 4709 3924 4721 3927
rect 4672 3896 4721 3924
rect 4672 3884 4678 3896
rect 4709 3893 4721 3896
rect 4755 3893 4767 3927
rect 4709 3887 4767 3893
rect 5350 3884 5356 3936
rect 5408 3884 5414 3936
rect 1104 3834 5796 3856
rect 1104 3782 1950 3834
rect 2002 3782 2014 3834
rect 2066 3782 2078 3834
rect 2130 3782 2142 3834
rect 2194 3782 2206 3834
rect 2258 3782 5796 3834
rect 1104 3760 5796 3782
rect 3234 3544 3240 3596
rect 3292 3584 3298 3596
rect 4617 3587 4675 3593
rect 4617 3584 4629 3587
rect 3292 3556 4629 3584
rect 3292 3544 3298 3556
rect 4617 3553 4629 3556
rect 4663 3553 4675 3587
rect 4617 3547 4675 3553
rect 5074 3544 5080 3596
rect 5132 3544 5138 3596
rect 4706 3476 4712 3528
rect 4764 3476 4770 3528
rect 1104 3290 5796 3312
rect 1104 3238 2610 3290
rect 2662 3238 2674 3290
rect 2726 3238 2738 3290
rect 2790 3238 2802 3290
rect 2854 3238 2866 3290
rect 2918 3238 5796 3290
rect 1104 3216 5796 3238
rect 4798 3136 4804 3188
rect 4856 3176 4862 3188
rect 4893 3179 4951 3185
rect 4893 3176 4905 3179
rect 4856 3148 4905 3176
rect 4856 3136 4862 3148
rect 4893 3145 4905 3148
rect 4939 3145 4951 3179
rect 4893 3139 4951 3145
rect 4341 3111 4399 3117
rect 4341 3077 4353 3111
rect 4387 3108 4399 3111
rect 4982 3108 4988 3120
rect 4387 3080 4988 3108
rect 4387 3077 4399 3080
rect 4341 3071 4399 3077
rect 4982 3068 4988 3080
rect 5040 3068 5046 3120
rect 4246 3000 4252 3052
rect 4304 3000 4310 3052
rect 4430 3000 4436 3052
rect 4488 3000 4494 3052
rect 5077 3043 5135 3049
rect 5077 3009 5089 3043
rect 5123 3009 5135 3043
rect 5077 3003 5135 3009
rect 3970 2932 3976 2984
rect 4028 2972 4034 2984
rect 5092 2972 5120 3003
rect 5258 3000 5264 3052
rect 5316 3000 5322 3052
rect 5353 3043 5411 3049
rect 5353 3009 5365 3043
rect 5399 3040 5411 3043
rect 5442 3040 5448 3052
rect 5399 3012 5448 3040
rect 5399 3009 5411 3012
rect 5353 3003 5411 3009
rect 5442 3000 5448 3012
rect 5500 3000 5506 3052
rect 4028 2944 5120 2972
rect 4028 2932 4034 2944
rect 3786 2864 3792 2916
rect 3844 2904 3850 2916
rect 5169 2907 5227 2913
rect 5169 2904 5181 2907
rect 3844 2876 5181 2904
rect 3844 2864 3850 2876
rect 5169 2873 5181 2876
rect 5215 2873 5227 2907
rect 5169 2867 5227 2873
rect 1104 2746 5796 2768
rect 1104 2694 1950 2746
rect 2002 2694 2014 2746
rect 2066 2694 2078 2746
rect 2130 2694 2142 2746
rect 2194 2694 2206 2746
rect 2258 2694 5796 2746
rect 1104 2672 5796 2694
rect 1857 2635 1915 2641
rect 1857 2601 1869 2635
rect 1903 2632 1915 2635
rect 4706 2632 4712 2644
rect 1903 2604 4712 2632
rect 1903 2601 1915 2604
rect 1857 2595 1915 2601
rect 4706 2592 4712 2604
rect 4764 2592 4770 2644
rect 1581 2567 1639 2573
rect 1581 2533 1593 2567
rect 1627 2564 1639 2567
rect 2958 2564 2964 2576
rect 1627 2536 2964 2564
rect 1627 2533 1639 2536
rect 1581 2527 1639 2533
rect 2958 2524 2964 2536
rect 3016 2524 3022 2576
rect 4341 2567 4399 2573
rect 4341 2533 4353 2567
rect 4387 2564 4399 2567
rect 5166 2564 5172 2576
rect 4387 2536 5172 2564
rect 4387 2533 4399 2536
rect 4341 2527 4399 2533
rect 5166 2524 5172 2536
rect 5224 2524 5230 2576
rect 4065 2499 4123 2505
rect 4065 2465 4077 2499
rect 4111 2496 4123 2499
rect 4430 2496 4436 2508
rect 4111 2468 4436 2496
rect 4111 2465 4123 2468
rect 4065 2459 4123 2465
rect 4430 2456 4436 2468
rect 4488 2456 4494 2508
rect 842 2388 848 2440
rect 900 2428 906 2440
rect 1397 2431 1455 2437
rect 1397 2428 1409 2431
rect 900 2400 1409 2428
rect 900 2388 906 2400
rect 1397 2397 1409 2400
rect 1443 2397 1455 2431
rect 1397 2391 1455 2397
rect 1670 2388 1676 2440
rect 1728 2388 1734 2440
rect 3050 2388 3056 2440
rect 3108 2428 3114 2440
rect 3973 2431 4031 2437
rect 3973 2428 3985 2431
rect 3108 2400 3985 2428
rect 3108 2388 3114 2400
rect 3973 2397 3985 2400
rect 4019 2397 4031 2431
rect 3973 2391 4031 2397
rect 4614 2388 4620 2440
rect 4672 2388 4678 2440
rect 5074 2388 5080 2440
rect 5132 2388 5138 2440
rect 5442 2320 5448 2372
rect 5500 2320 5506 2372
rect 4798 2252 4804 2304
rect 4856 2252 4862 2304
rect 1104 2202 5796 2224
rect 1104 2150 2610 2202
rect 2662 2150 2674 2202
rect 2726 2150 2738 2202
rect 2790 2150 2802 2202
rect 2854 2150 2866 2202
rect 2918 2150 5796 2202
rect 1104 2128 5796 2150
<< via1 >>
rect 1950 9222 2002 9274
rect 2014 9222 2066 9274
rect 2078 9222 2130 9274
rect 2142 9222 2194 9274
rect 2206 9222 2258 9274
rect 4988 9163 5040 9172
rect 4988 9129 4997 9163
rect 4997 9129 5031 9163
rect 5031 9129 5040 9163
rect 4988 9120 5040 9129
rect 3056 9052 3108 9104
rect 5356 9095 5408 9104
rect 5356 9061 5365 9095
rect 5365 9061 5399 9095
rect 5399 9061 5408 9095
rect 5356 9052 5408 9061
rect 1400 8959 1452 8968
rect 1400 8925 1409 8959
rect 1409 8925 1443 8959
rect 1443 8925 1452 8959
rect 1400 8916 1452 8925
rect 3424 8984 3476 9036
rect 848 8848 900 8900
rect 3148 8916 3200 8968
rect 3516 8916 3568 8968
rect 5172 8959 5224 8968
rect 5172 8925 5181 8959
rect 5181 8925 5215 8959
rect 5215 8925 5224 8959
rect 5172 8916 5224 8925
rect 4344 8848 4396 8900
rect 1584 8823 1636 8832
rect 1584 8789 1593 8823
rect 1593 8789 1627 8823
rect 1627 8789 1636 8823
rect 1584 8780 1636 8789
rect 2964 8780 3016 8832
rect 3976 8780 4028 8832
rect 2610 8678 2662 8730
rect 2674 8678 2726 8730
rect 2738 8678 2790 8730
rect 2802 8678 2854 8730
rect 2866 8678 2918 8730
rect 3516 8619 3568 8628
rect 3516 8585 3525 8619
rect 3525 8585 3559 8619
rect 3559 8585 3568 8619
rect 3516 8576 3568 8585
rect 2412 8440 2464 8492
rect 2964 8483 3016 8492
rect 2964 8449 2973 8483
rect 2973 8449 3007 8483
rect 3007 8449 3016 8483
rect 2964 8440 3016 8449
rect 3332 8483 3384 8492
rect 2780 8415 2832 8424
rect 2780 8381 2789 8415
rect 2789 8381 2823 8415
rect 2823 8381 2832 8415
rect 2780 8372 2832 8381
rect 1584 8304 1636 8356
rect 3332 8449 3341 8483
rect 3341 8449 3375 8483
rect 3375 8449 3384 8483
rect 3332 8440 3384 8449
rect 3424 8372 3476 8424
rect 4344 8440 4396 8492
rect 4068 8415 4120 8424
rect 4068 8381 4077 8415
rect 4077 8381 4111 8415
rect 4111 8381 4120 8415
rect 4068 8372 4120 8381
rect 4436 8304 4488 8356
rect 1950 8134 2002 8186
rect 2014 8134 2066 8186
rect 2078 8134 2130 8186
rect 2142 8134 2194 8186
rect 2206 8134 2258 8186
rect 2504 8032 2556 8084
rect 2780 8032 2832 8084
rect 5172 7964 5224 8016
rect 1584 7871 1636 7880
rect 1584 7837 1593 7871
rect 1593 7837 1627 7871
rect 1627 7837 1636 7871
rect 1584 7828 1636 7837
rect 1768 7871 1820 7880
rect 1768 7837 1777 7871
rect 1777 7837 1811 7871
rect 1811 7837 1820 7871
rect 1768 7828 1820 7837
rect 940 7760 992 7812
rect 4160 7828 4212 7880
rect 5356 7735 5408 7744
rect 5356 7701 5365 7735
rect 5365 7701 5399 7735
rect 5399 7701 5408 7735
rect 5356 7692 5408 7701
rect 2610 7590 2662 7642
rect 2674 7590 2726 7642
rect 2738 7590 2790 7642
rect 2802 7590 2854 7642
rect 2866 7590 2918 7642
rect 1768 7488 1820 7540
rect 2964 7420 3016 7472
rect 3332 7395 3384 7404
rect 3332 7361 3341 7395
rect 3341 7361 3375 7395
rect 3375 7361 3384 7395
rect 3332 7352 3384 7361
rect 3884 7420 3936 7472
rect 3976 7352 4028 7404
rect 3792 7284 3844 7336
rect 3240 7216 3292 7268
rect 4252 7191 4304 7200
rect 4252 7157 4261 7191
rect 4261 7157 4295 7191
rect 4295 7157 4304 7191
rect 4252 7148 4304 7157
rect 1950 7046 2002 7098
rect 2014 7046 2066 7098
rect 2078 7046 2130 7098
rect 2142 7046 2194 7098
rect 2206 7046 2258 7098
rect 4344 6808 4396 6860
rect 848 6740 900 6792
rect 2412 6604 2464 6656
rect 5448 6740 5500 6792
rect 4804 6715 4856 6724
rect 4804 6681 4813 6715
rect 4813 6681 4847 6715
rect 4847 6681 4856 6715
rect 4804 6672 4856 6681
rect 4896 6604 4948 6656
rect 2610 6502 2662 6554
rect 2674 6502 2726 6554
rect 2738 6502 2790 6554
rect 2802 6502 2854 6554
rect 2866 6502 2918 6554
rect 5356 6443 5408 6452
rect 5356 6409 5365 6443
rect 5365 6409 5399 6443
rect 5399 6409 5408 6443
rect 5356 6400 5408 6409
rect 5172 6307 5224 6316
rect 5172 6273 5181 6307
rect 5181 6273 5215 6307
rect 5215 6273 5224 6307
rect 5172 6264 5224 6273
rect 1950 5958 2002 6010
rect 2014 5958 2066 6010
rect 2078 5958 2130 6010
rect 2142 5958 2194 6010
rect 2206 5958 2258 6010
rect 4160 5788 4212 5840
rect 1584 5720 1636 5772
rect 2504 5695 2556 5704
rect 2504 5661 2513 5695
rect 2513 5661 2547 5695
rect 2547 5661 2556 5695
rect 2504 5652 2556 5661
rect 3792 5695 3844 5704
rect 3792 5661 3801 5695
rect 3801 5661 3835 5695
rect 3835 5661 3844 5695
rect 3792 5652 3844 5661
rect 3976 5695 4028 5704
rect 3976 5661 3985 5695
rect 3985 5661 4019 5695
rect 4019 5661 4028 5695
rect 3976 5652 4028 5661
rect 5264 5584 5316 5636
rect 2610 5414 2662 5466
rect 2674 5414 2726 5466
rect 2738 5414 2790 5466
rect 2802 5414 2854 5466
rect 2866 5414 2918 5466
rect 848 5176 900 5228
rect 5172 5312 5224 5364
rect 3332 5176 3384 5228
rect 4896 5219 4948 5228
rect 4896 5185 4905 5219
rect 4905 5185 4939 5219
rect 4939 5185 4948 5219
rect 4896 5176 4948 5185
rect 4988 5176 5040 5228
rect 2964 5151 3016 5160
rect 2964 5117 2973 5151
rect 2973 5117 3007 5151
rect 3007 5117 3016 5151
rect 2964 5108 3016 5117
rect 3148 5108 3200 5160
rect 4344 5040 4396 5092
rect 3056 5015 3108 5024
rect 3056 4981 3065 5015
rect 3065 4981 3099 5015
rect 3099 4981 3108 5015
rect 3056 4972 3108 4981
rect 3240 5015 3292 5024
rect 3240 4981 3249 5015
rect 3249 4981 3283 5015
rect 3283 4981 3292 5015
rect 3240 4972 3292 4981
rect 5356 5015 5408 5024
rect 5356 4981 5365 5015
rect 5365 4981 5399 5015
rect 5399 4981 5408 5015
rect 5356 4972 5408 4981
rect 1950 4870 2002 4922
rect 2014 4870 2066 4922
rect 2078 4870 2130 4922
rect 2142 4870 2194 4922
rect 2206 4870 2258 4922
rect 2610 4326 2662 4378
rect 2674 4326 2726 4378
rect 2738 4326 2790 4378
rect 2802 4326 2854 4378
rect 2866 4326 2918 4378
rect 848 4088 900 4140
rect 4252 4088 4304 4140
rect 5172 4131 5224 4140
rect 5172 4097 5181 4131
rect 5181 4097 5215 4131
rect 5215 4097 5224 4131
rect 5172 4088 5224 4097
rect 3056 3952 3108 4004
rect 4620 3884 4672 3936
rect 5356 3927 5408 3936
rect 5356 3893 5365 3927
rect 5365 3893 5399 3927
rect 5399 3893 5408 3927
rect 5356 3884 5408 3893
rect 1950 3782 2002 3834
rect 2014 3782 2066 3834
rect 2078 3782 2130 3834
rect 2142 3782 2194 3834
rect 2206 3782 2258 3834
rect 3240 3544 3292 3596
rect 5080 3587 5132 3596
rect 5080 3553 5089 3587
rect 5089 3553 5123 3587
rect 5123 3553 5132 3587
rect 5080 3544 5132 3553
rect 4712 3519 4764 3528
rect 4712 3485 4721 3519
rect 4721 3485 4755 3519
rect 4755 3485 4764 3519
rect 4712 3476 4764 3485
rect 2610 3238 2662 3290
rect 2674 3238 2726 3290
rect 2738 3238 2790 3290
rect 2802 3238 2854 3290
rect 2866 3238 2918 3290
rect 4804 3136 4856 3188
rect 4988 3068 5040 3120
rect 4252 3043 4304 3052
rect 4252 3009 4261 3043
rect 4261 3009 4295 3043
rect 4295 3009 4304 3043
rect 4252 3000 4304 3009
rect 4436 3043 4488 3052
rect 4436 3009 4445 3043
rect 4445 3009 4479 3043
rect 4479 3009 4488 3043
rect 4436 3000 4488 3009
rect 3976 2932 4028 2984
rect 5264 3043 5316 3052
rect 5264 3009 5273 3043
rect 5273 3009 5307 3043
rect 5307 3009 5316 3043
rect 5264 3000 5316 3009
rect 5448 3000 5500 3052
rect 3792 2864 3844 2916
rect 1950 2694 2002 2746
rect 2014 2694 2066 2746
rect 2078 2694 2130 2746
rect 2142 2694 2194 2746
rect 2206 2694 2258 2746
rect 4712 2592 4764 2644
rect 2964 2524 3016 2576
rect 5172 2524 5224 2576
rect 4436 2456 4488 2508
rect 848 2388 900 2440
rect 1676 2431 1728 2440
rect 1676 2397 1685 2431
rect 1685 2397 1719 2431
rect 1719 2397 1728 2431
rect 1676 2388 1728 2397
rect 3056 2388 3108 2440
rect 4620 2431 4672 2440
rect 4620 2397 4629 2431
rect 4629 2397 4663 2431
rect 4663 2397 4672 2431
rect 4620 2388 4672 2397
rect 5080 2431 5132 2440
rect 5080 2397 5089 2431
rect 5089 2397 5123 2431
rect 5123 2397 5132 2431
rect 5080 2388 5132 2397
rect 5448 2363 5500 2372
rect 5448 2329 5457 2363
rect 5457 2329 5491 2363
rect 5491 2329 5500 2363
rect 5448 2320 5500 2329
rect 4804 2295 4856 2304
rect 4804 2261 4813 2295
rect 4813 2261 4847 2295
rect 4847 2261 4856 2295
rect 4804 2252 4856 2261
rect 2610 2150 2662 2202
rect 2674 2150 2726 2202
rect 2738 2150 2790 2202
rect 2802 2150 2854 2202
rect 2866 2150 2918 2202
<< metal2 >>
rect 1398 10432 1454 10441
rect 1398 10367 1454 10376
rect 4986 10432 5042 10441
rect 4986 10367 5042 10376
rect 1412 8974 1440 10367
rect 1950 9276 2258 9285
rect 1950 9274 1956 9276
rect 2012 9274 2036 9276
rect 2092 9274 2116 9276
rect 2172 9274 2196 9276
rect 2252 9274 2258 9276
rect 2012 9222 2014 9274
rect 2194 9222 2196 9274
rect 1950 9220 1956 9222
rect 2012 9220 2036 9222
rect 2092 9220 2116 9222
rect 2172 9220 2196 9222
rect 2252 9220 2258 9222
rect 1950 9211 2258 9220
rect 5000 9178 5028 10367
rect 4988 9172 5040 9178
rect 4988 9114 5040 9120
rect 3056 9104 3108 9110
rect 5356 9104 5408 9110
rect 3056 9046 3108 9052
rect 5354 9072 5356 9081
rect 5408 9072 5410 9081
rect 1400 8968 1452 8974
rect 846 8936 902 8945
rect 1400 8910 1452 8916
rect 846 8871 848 8880
rect 900 8871 902 8880
rect 848 8842 900 8848
rect 1584 8832 1636 8838
rect 1584 8774 1636 8780
rect 2964 8832 3016 8838
rect 2964 8774 3016 8780
rect 1596 8362 1624 8774
rect 2610 8732 2918 8741
rect 2610 8730 2616 8732
rect 2672 8730 2696 8732
rect 2752 8730 2776 8732
rect 2832 8730 2856 8732
rect 2912 8730 2918 8732
rect 2672 8678 2674 8730
rect 2854 8678 2856 8730
rect 2610 8676 2616 8678
rect 2672 8676 2696 8678
rect 2752 8676 2776 8678
rect 2832 8676 2856 8678
rect 2912 8676 2918 8678
rect 2610 8667 2918 8676
rect 2976 8498 3004 8774
rect 2412 8492 2464 8498
rect 2412 8434 2464 8440
rect 2964 8492 3016 8498
rect 2964 8434 3016 8440
rect 1584 8356 1636 8362
rect 1584 8298 1636 8304
rect 1950 8188 2258 8197
rect 1950 8186 1956 8188
rect 2012 8186 2036 8188
rect 2092 8186 2116 8188
rect 2172 8186 2196 8188
rect 2252 8186 2258 8188
rect 2012 8134 2014 8186
rect 2194 8134 2196 8186
rect 1950 8132 1956 8134
rect 2012 8132 2036 8134
rect 2092 8132 2116 8134
rect 2172 8132 2196 8134
rect 2252 8132 2258 8134
rect 1950 8123 2258 8132
rect 1584 7880 1636 7886
rect 1584 7822 1636 7828
rect 1768 7880 1820 7886
rect 1768 7822 1820 7828
rect 940 7812 992 7818
rect 940 7754 992 7760
rect 952 7721 980 7754
rect 938 7712 994 7721
rect 938 7647 994 7656
rect 848 6792 900 6798
rect 848 6734 900 6740
rect 860 6497 888 6734
rect 846 6488 902 6497
rect 846 6423 902 6432
rect 1596 5778 1624 7822
rect 1780 7546 1808 7822
rect 1768 7540 1820 7546
rect 1768 7482 1820 7488
rect 1950 7100 2258 7109
rect 1950 7098 1956 7100
rect 2012 7098 2036 7100
rect 2092 7098 2116 7100
rect 2172 7098 2196 7100
rect 2252 7098 2258 7100
rect 2012 7046 2014 7098
rect 2194 7046 2196 7098
rect 1950 7044 1956 7046
rect 2012 7044 2036 7046
rect 2092 7044 2116 7046
rect 2172 7044 2196 7046
rect 2252 7044 2258 7046
rect 1950 7035 2258 7044
rect 2424 6662 2452 8434
rect 2780 8424 2832 8430
rect 2780 8366 2832 8372
rect 2792 8090 2820 8366
rect 2504 8084 2556 8090
rect 2504 8026 2556 8032
rect 2780 8084 2832 8090
rect 2780 8026 2832 8032
rect 2412 6656 2464 6662
rect 2412 6598 2464 6604
rect 1950 6012 2258 6021
rect 1950 6010 1956 6012
rect 2012 6010 2036 6012
rect 2092 6010 2116 6012
rect 2172 6010 2196 6012
rect 2252 6010 2258 6012
rect 2012 5958 2014 6010
rect 2194 5958 2196 6010
rect 1950 5956 1956 5958
rect 2012 5956 2036 5958
rect 2092 5956 2116 5958
rect 2172 5956 2196 5958
rect 2252 5956 2258 5958
rect 1950 5947 2258 5956
rect 1584 5772 1636 5778
rect 1584 5714 1636 5720
rect 2516 5710 2544 8026
rect 2610 7644 2918 7653
rect 2610 7642 2616 7644
rect 2672 7642 2696 7644
rect 2752 7642 2776 7644
rect 2832 7642 2856 7644
rect 2912 7642 2918 7644
rect 2672 7590 2674 7642
rect 2854 7590 2856 7642
rect 2610 7588 2616 7590
rect 2672 7588 2696 7590
rect 2752 7588 2776 7590
rect 2832 7588 2856 7590
rect 2912 7588 2918 7590
rect 2610 7579 2918 7588
rect 2976 7478 3004 8434
rect 2964 7472 3016 7478
rect 2964 7414 3016 7420
rect 2610 6556 2918 6565
rect 2610 6554 2616 6556
rect 2672 6554 2696 6556
rect 2752 6554 2776 6556
rect 2832 6554 2856 6556
rect 2912 6554 2918 6556
rect 2672 6502 2674 6554
rect 2854 6502 2856 6554
rect 2610 6500 2616 6502
rect 2672 6500 2696 6502
rect 2752 6500 2776 6502
rect 2832 6500 2856 6502
rect 2912 6500 2918 6502
rect 2610 6491 2918 6500
rect 2504 5704 2556 5710
rect 2504 5646 2556 5652
rect 2610 5468 2918 5477
rect 2610 5466 2616 5468
rect 2672 5466 2696 5468
rect 2752 5466 2776 5468
rect 2832 5466 2856 5468
rect 2912 5466 2918 5468
rect 2672 5414 2674 5466
rect 2854 5414 2856 5466
rect 2610 5412 2616 5414
rect 2672 5412 2696 5414
rect 2752 5412 2776 5414
rect 2832 5412 2856 5414
rect 2912 5412 2918 5414
rect 2610 5403 2918 5412
rect 848 5228 900 5234
rect 848 5170 900 5176
rect 860 5137 888 5170
rect 2964 5160 3016 5166
rect 846 5128 902 5137
rect 2964 5102 3016 5108
rect 846 5063 902 5072
rect 1950 4924 2258 4933
rect 1950 4922 1956 4924
rect 2012 4922 2036 4924
rect 2092 4922 2116 4924
rect 2172 4922 2196 4924
rect 2252 4922 2258 4924
rect 2012 4870 2014 4922
rect 2194 4870 2196 4922
rect 1950 4868 1956 4870
rect 2012 4868 2036 4870
rect 2092 4868 2116 4870
rect 2172 4868 2196 4870
rect 2252 4868 2258 4870
rect 1950 4859 2258 4868
rect 2610 4380 2918 4389
rect 2610 4378 2616 4380
rect 2672 4378 2696 4380
rect 2752 4378 2776 4380
rect 2832 4378 2856 4380
rect 2912 4378 2918 4380
rect 2672 4326 2674 4378
rect 2854 4326 2856 4378
rect 2610 4324 2616 4326
rect 2672 4324 2696 4326
rect 2752 4324 2776 4326
rect 2832 4324 2856 4326
rect 2912 4324 2918 4326
rect 2610 4315 2918 4324
rect 848 4140 900 4146
rect 848 4082 900 4088
rect 860 3777 888 4082
rect 1950 3836 2258 3845
rect 1950 3834 1956 3836
rect 2012 3834 2036 3836
rect 2092 3834 2116 3836
rect 2172 3834 2196 3836
rect 2252 3834 2258 3836
rect 2012 3782 2014 3834
rect 2194 3782 2196 3834
rect 1950 3780 1956 3782
rect 2012 3780 2036 3782
rect 2092 3780 2116 3782
rect 2172 3780 2196 3782
rect 2252 3780 2258 3782
rect 846 3768 902 3777
rect 1950 3771 2258 3780
rect 846 3703 902 3712
rect 2610 3292 2918 3301
rect 2610 3290 2616 3292
rect 2672 3290 2696 3292
rect 2752 3290 2776 3292
rect 2832 3290 2856 3292
rect 2912 3290 2918 3292
rect 2672 3238 2674 3290
rect 2854 3238 2856 3290
rect 2610 3236 2616 3238
rect 2672 3236 2696 3238
rect 2752 3236 2776 3238
rect 2832 3236 2856 3238
rect 2912 3236 2918 3238
rect 2610 3227 2918 3236
rect 1950 2748 2258 2757
rect 1950 2746 1956 2748
rect 2012 2746 2036 2748
rect 2092 2746 2116 2748
rect 2172 2746 2196 2748
rect 2252 2746 2258 2748
rect 2012 2694 2014 2746
rect 2194 2694 2196 2746
rect 1950 2692 1956 2694
rect 2012 2692 2036 2694
rect 2092 2692 2116 2694
rect 2172 2692 2196 2694
rect 2252 2692 2258 2694
rect 1950 2683 2258 2692
rect 2976 2582 3004 5102
rect 3068 5030 3096 9046
rect 3424 9036 3476 9042
rect 5354 9007 5410 9016
rect 3424 8978 3476 8984
rect 3148 8968 3200 8974
rect 3148 8910 3200 8916
rect 3160 5166 3188 8910
rect 3332 8492 3384 8498
rect 3332 8434 3384 8440
rect 3344 7410 3372 8434
rect 3436 8430 3464 8978
rect 3516 8968 3568 8974
rect 3516 8910 3568 8916
rect 5172 8968 5224 8974
rect 5172 8910 5224 8916
rect 3528 8634 3556 8910
rect 4344 8900 4396 8906
rect 4344 8842 4396 8848
rect 3976 8832 4028 8838
rect 3976 8774 4028 8780
rect 3516 8628 3568 8634
rect 3516 8570 3568 8576
rect 3424 8424 3476 8430
rect 3424 8366 3476 8372
rect 3332 7404 3384 7410
rect 3332 7346 3384 7352
rect 3240 7268 3292 7274
rect 3240 7210 3292 7216
rect 3148 5160 3200 5166
rect 3148 5102 3200 5108
rect 3252 5030 3280 7210
rect 3436 6914 3464 8366
rect 3884 7472 3936 7478
rect 3884 7414 3936 7420
rect 3792 7336 3844 7342
rect 3792 7278 3844 7284
rect 3344 6886 3464 6914
rect 3344 5234 3372 6886
rect 3804 5710 3832 7278
rect 3896 6914 3924 7414
rect 3988 7410 4016 8774
rect 4356 8498 4384 8842
rect 4344 8492 4396 8498
rect 4344 8434 4396 8440
rect 4068 8424 4120 8430
rect 4066 8392 4068 8401
rect 4120 8392 4122 8401
rect 4066 8327 4122 8336
rect 4160 7880 4212 7886
rect 4160 7822 4212 7828
rect 3976 7404 4028 7410
rect 3976 7346 4028 7352
rect 3896 6886 4016 6914
rect 3988 5710 4016 6886
rect 4172 5846 4200 7822
rect 4252 7200 4304 7206
rect 4252 7142 4304 7148
rect 4160 5840 4212 5846
rect 4160 5782 4212 5788
rect 3792 5704 3844 5710
rect 3792 5646 3844 5652
rect 3976 5704 4028 5710
rect 3976 5646 4028 5652
rect 3332 5228 3384 5234
rect 3332 5170 3384 5176
rect 3056 5024 3108 5030
rect 3056 4966 3108 4972
rect 3240 5024 3292 5030
rect 3240 4966 3292 4972
rect 3068 4010 3096 4966
rect 3056 4004 3108 4010
rect 3056 3946 3108 3952
rect 2964 2576 3016 2582
rect 2964 2518 3016 2524
rect 3068 2446 3096 3946
rect 3252 3602 3280 4966
rect 3240 3596 3292 3602
rect 3240 3538 3292 3544
rect 3804 2922 3832 5646
rect 3988 2990 4016 5646
rect 4264 4146 4292 7142
rect 4356 6866 4384 8434
rect 4436 8356 4488 8362
rect 4436 8298 4488 8304
rect 4344 6860 4396 6866
rect 4344 6802 4396 6808
rect 4356 5098 4384 6802
rect 4344 5092 4396 5098
rect 4344 5034 4396 5040
rect 4252 4140 4304 4146
rect 4252 4082 4304 4088
rect 4250 4040 4306 4049
rect 4250 3975 4306 3984
rect 4264 3058 4292 3975
rect 4448 3058 4476 8298
rect 5184 8022 5212 8910
rect 5172 8016 5224 8022
rect 5172 7958 5224 7964
rect 5356 7744 5408 7750
rect 5354 7712 5356 7721
rect 5408 7712 5410 7721
rect 5354 7647 5410 7656
rect 5448 6792 5500 6798
rect 5448 6734 5500 6740
rect 4804 6724 4856 6730
rect 4804 6666 4856 6672
rect 4620 3936 4672 3942
rect 4620 3878 4672 3884
rect 4252 3052 4304 3058
rect 4252 2994 4304 3000
rect 4436 3052 4488 3058
rect 4436 2994 4488 3000
rect 3976 2984 4028 2990
rect 3976 2926 4028 2932
rect 3792 2916 3844 2922
rect 3792 2858 3844 2864
rect 4448 2514 4476 2994
rect 4436 2508 4488 2514
rect 4436 2450 4488 2456
rect 4632 2446 4660 3878
rect 4712 3528 4764 3534
rect 4712 3470 4764 3476
rect 4724 2650 4752 3470
rect 4816 3194 4844 6666
rect 4896 6656 4948 6662
rect 4896 6598 4948 6604
rect 4908 5234 4936 6598
rect 5356 6452 5408 6458
rect 5356 6394 5408 6400
rect 5368 6361 5396 6394
rect 5354 6352 5410 6361
rect 5172 6316 5224 6322
rect 5354 6287 5410 6296
rect 5172 6258 5224 6264
rect 5184 5370 5212 6258
rect 5264 5636 5316 5642
rect 5264 5578 5316 5584
rect 5172 5364 5224 5370
rect 5172 5306 5224 5312
rect 4896 5228 4948 5234
rect 4896 5170 4948 5176
rect 4988 5228 5040 5234
rect 4988 5170 5040 5176
rect 4804 3188 4856 3194
rect 4804 3130 4856 3136
rect 5000 3126 5028 5170
rect 5172 4140 5224 4146
rect 5172 4082 5224 4088
rect 5080 3596 5132 3602
rect 5080 3538 5132 3544
rect 4988 3120 5040 3126
rect 4988 3062 5040 3068
rect 4712 2644 4764 2650
rect 4712 2586 4764 2592
rect 5092 2446 5120 3538
rect 5184 2582 5212 4082
rect 5276 3058 5304 5578
rect 5356 5024 5408 5030
rect 5354 4992 5356 5001
rect 5408 4992 5410 5001
rect 5354 4927 5410 4936
rect 5356 3936 5408 3942
rect 5356 3878 5408 3884
rect 5368 3641 5396 3878
rect 5354 3632 5410 3641
rect 5354 3567 5410 3576
rect 5460 3058 5488 6734
rect 5264 3052 5316 3058
rect 5264 2994 5316 3000
rect 5448 3052 5500 3058
rect 5448 2994 5500 3000
rect 5172 2576 5224 2582
rect 5172 2518 5224 2524
rect 848 2440 900 2446
rect 846 2408 848 2417
rect 1676 2440 1728 2446
rect 900 2408 902 2417
rect 1676 2382 1728 2388
rect 3056 2440 3108 2446
rect 3056 2382 3108 2388
rect 4620 2440 4672 2446
rect 4620 2382 4672 2388
rect 5080 2440 5132 2446
rect 5080 2382 5132 2388
rect 846 2343 902 2352
rect 1688 921 1716 2382
rect 5448 2372 5500 2378
rect 5448 2314 5500 2320
rect 4804 2304 4856 2310
rect 4802 2272 4804 2281
rect 4856 2272 4858 2281
rect 2610 2204 2918 2213
rect 4802 2207 4858 2216
rect 2610 2202 2616 2204
rect 2672 2202 2696 2204
rect 2752 2202 2776 2204
rect 2832 2202 2856 2204
rect 2912 2202 2918 2204
rect 2672 2150 2674 2202
rect 2854 2150 2856 2202
rect 2610 2148 2616 2150
rect 2672 2148 2696 2150
rect 2752 2148 2776 2150
rect 2832 2148 2856 2150
rect 2912 2148 2918 2150
rect 2610 2139 2918 2148
rect 5460 921 5488 2314
rect 1674 912 1730 921
rect 1674 847 1730 856
rect 5446 912 5502 921
rect 5446 847 5502 856
<< via2 >>
rect 1398 10376 1454 10432
rect 4986 10376 5042 10432
rect 1956 9274 2012 9276
rect 2036 9274 2092 9276
rect 2116 9274 2172 9276
rect 2196 9274 2252 9276
rect 1956 9222 2002 9274
rect 2002 9222 2012 9274
rect 2036 9222 2066 9274
rect 2066 9222 2078 9274
rect 2078 9222 2092 9274
rect 2116 9222 2130 9274
rect 2130 9222 2142 9274
rect 2142 9222 2172 9274
rect 2196 9222 2206 9274
rect 2206 9222 2252 9274
rect 1956 9220 2012 9222
rect 2036 9220 2092 9222
rect 2116 9220 2172 9222
rect 2196 9220 2252 9222
rect 5354 9052 5356 9072
rect 5356 9052 5408 9072
rect 5408 9052 5410 9072
rect 846 8900 902 8936
rect 846 8880 848 8900
rect 848 8880 900 8900
rect 900 8880 902 8900
rect 2616 8730 2672 8732
rect 2696 8730 2752 8732
rect 2776 8730 2832 8732
rect 2856 8730 2912 8732
rect 2616 8678 2662 8730
rect 2662 8678 2672 8730
rect 2696 8678 2726 8730
rect 2726 8678 2738 8730
rect 2738 8678 2752 8730
rect 2776 8678 2790 8730
rect 2790 8678 2802 8730
rect 2802 8678 2832 8730
rect 2856 8678 2866 8730
rect 2866 8678 2912 8730
rect 2616 8676 2672 8678
rect 2696 8676 2752 8678
rect 2776 8676 2832 8678
rect 2856 8676 2912 8678
rect 1956 8186 2012 8188
rect 2036 8186 2092 8188
rect 2116 8186 2172 8188
rect 2196 8186 2252 8188
rect 1956 8134 2002 8186
rect 2002 8134 2012 8186
rect 2036 8134 2066 8186
rect 2066 8134 2078 8186
rect 2078 8134 2092 8186
rect 2116 8134 2130 8186
rect 2130 8134 2142 8186
rect 2142 8134 2172 8186
rect 2196 8134 2206 8186
rect 2206 8134 2252 8186
rect 1956 8132 2012 8134
rect 2036 8132 2092 8134
rect 2116 8132 2172 8134
rect 2196 8132 2252 8134
rect 938 7656 994 7712
rect 846 6432 902 6488
rect 1956 7098 2012 7100
rect 2036 7098 2092 7100
rect 2116 7098 2172 7100
rect 2196 7098 2252 7100
rect 1956 7046 2002 7098
rect 2002 7046 2012 7098
rect 2036 7046 2066 7098
rect 2066 7046 2078 7098
rect 2078 7046 2092 7098
rect 2116 7046 2130 7098
rect 2130 7046 2142 7098
rect 2142 7046 2172 7098
rect 2196 7046 2206 7098
rect 2206 7046 2252 7098
rect 1956 7044 2012 7046
rect 2036 7044 2092 7046
rect 2116 7044 2172 7046
rect 2196 7044 2252 7046
rect 1956 6010 2012 6012
rect 2036 6010 2092 6012
rect 2116 6010 2172 6012
rect 2196 6010 2252 6012
rect 1956 5958 2002 6010
rect 2002 5958 2012 6010
rect 2036 5958 2066 6010
rect 2066 5958 2078 6010
rect 2078 5958 2092 6010
rect 2116 5958 2130 6010
rect 2130 5958 2142 6010
rect 2142 5958 2172 6010
rect 2196 5958 2206 6010
rect 2206 5958 2252 6010
rect 1956 5956 2012 5958
rect 2036 5956 2092 5958
rect 2116 5956 2172 5958
rect 2196 5956 2252 5958
rect 2616 7642 2672 7644
rect 2696 7642 2752 7644
rect 2776 7642 2832 7644
rect 2856 7642 2912 7644
rect 2616 7590 2662 7642
rect 2662 7590 2672 7642
rect 2696 7590 2726 7642
rect 2726 7590 2738 7642
rect 2738 7590 2752 7642
rect 2776 7590 2790 7642
rect 2790 7590 2802 7642
rect 2802 7590 2832 7642
rect 2856 7590 2866 7642
rect 2866 7590 2912 7642
rect 2616 7588 2672 7590
rect 2696 7588 2752 7590
rect 2776 7588 2832 7590
rect 2856 7588 2912 7590
rect 2616 6554 2672 6556
rect 2696 6554 2752 6556
rect 2776 6554 2832 6556
rect 2856 6554 2912 6556
rect 2616 6502 2662 6554
rect 2662 6502 2672 6554
rect 2696 6502 2726 6554
rect 2726 6502 2738 6554
rect 2738 6502 2752 6554
rect 2776 6502 2790 6554
rect 2790 6502 2802 6554
rect 2802 6502 2832 6554
rect 2856 6502 2866 6554
rect 2866 6502 2912 6554
rect 2616 6500 2672 6502
rect 2696 6500 2752 6502
rect 2776 6500 2832 6502
rect 2856 6500 2912 6502
rect 2616 5466 2672 5468
rect 2696 5466 2752 5468
rect 2776 5466 2832 5468
rect 2856 5466 2912 5468
rect 2616 5414 2662 5466
rect 2662 5414 2672 5466
rect 2696 5414 2726 5466
rect 2726 5414 2738 5466
rect 2738 5414 2752 5466
rect 2776 5414 2790 5466
rect 2790 5414 2802 5466
rect 2802 5414 2832 5466
rect 2856 5414 2866 5466
rect 2866 5414 2912 5466
rect 2616 5412 2672 5414
rect 2696 5412 2752 5414
rect 2776 5412 2832 5414
rect 2856 5412 2912 5414
rect 846 5072 902 5128
rect 1956 4922 2012 4924
rect 2036 4922 2092 4924
rect 2116 4922 2172 4924
rect 2196 4922 2252 4924
rect 1956 4870 2002 4922
rect 2002 4870 2012 4922
rect 2036 4870 2066 4922
rect 2066 4870 2078 4922
rect 2078 4870 2092 4922
rect 2116 4870 2130 4922
rect 2130 4870 2142 4922
rect 2142 4870 2172 4922
rect 2196 4870 2206 4922
rect 2206 4870 2252 4922
rect 1956 4868 2012 4870
rect 2036 4868 2092 4870
rect 2116 4868 2172 4870
rect 2196 4868 2252 4870
rect 2616 4378 2672 4380
rect 2696 4378 2752 4380
rect 2776 4378 2832 4380
rect 2856 4378 2912 4380
rect 2616 4326 2662 4378
rect 2662 4326 2672 4378
rect 2696 4326 2726 4378
rect 2726 4326 2738 4378
rect 2738 4326 2752 4378
rect 2776 4326 2790 4378
rect 2790 4326 2802 4378
rect 2802 4326 2832 4378
rect 2856 4326 2866 4378
rect 2866 4326 2912 4378
rect 2616 4324 2672 4326
rect 2696 4324 2752 4326
rect 2776 4324 2832 4326
rect 2856 4324 2912 4326
rect 1956 3834 2012 3836
rect 2036 3834 2092 3836
rect 2116 3834 2172 3836
rect 2196 3834 2252 3836
rect 1956 3782 2002 3834
rect 2002 3782 2012 3834
rect 2036 3782 2066 3834
rect 2066 3782 2078 3834
rect 2078 3782 2092 3834
rect 2116 3782 2130 3834
rect 2130 3782 2142 3834
rect 2142 3782 2172 3834
rect 2196 3782 2206 3834
rect 2206 3782 2252 3834
rect 1956 3780 2012 3782
rect 2036 3780 2092 3782
rect 2116 3780 2172 3782
rect 2196 3780 2252 3782
rect 846 3712 902 3768
rect 2616 3290 2672 3292
rect 2696 3290 2752 3292
rect 2776 3290 2832 3292
rect 2856 3290 2912 3292
rect 2616 3238 2662 3290
rect 2662 3238 2672 3290
rect 2696 3238 2726 3290
rect 2726 3238 2738 3290
rect 2738 3238 2752 3290
rect 2776 3238 2790 3290
rect 2790 3238 2802 3290
rect 2802 3238 2832 3290
rect 2856 3238 2866 3290
rect 2866 3238 2912 3290
rect 2616 3236 2672 3238
rect 2696 3236 2752 3238
rect 2776 3236 2832 3238
rect 2856 3236 2912 3238
rect 1956 2746 2012 2748
rect 2036 2746 2092 2748
rect 2116 2746 2172 2748
rect 2196 2746 2252 2748
rect 1956 2694 2002 2746
rect 2002 2694 2012 2746
rect 2036 2694 2066 2746
rect 2066 2694 2078 2746
rect 2078 2694 2092 2746
rect 2116 2694 2130 2746
rect 2130 2694 2142 2746
rect 2142 2694 2172 2746
rect 2196 2694 2206 2746
rect 2206 2694 2252 2746
rect 1956 2692 2012 2694
rect 2036 2692 2092 2694
rect 2116 2692 2172 2694
rect 2196 2692 2252 2694
rect 5354 9016 5410 9052
rect 4066 8372 4068 8392
rect 4068 8372 4120 8392
rect 4120 8372 4122 8392
rect 4066 8336 4122 8372
rect 4250 3984 4306 4040
rect 5354 7692 5356 7712
rect 5356 7692 5408 7712
rect 5408 7692 5410 7712
rect 5354 7656 5410 7692
rect 5354 6296 5410 6352
rect 5354 4972 5356 4992
rect 5356 4972 5408 4992
rect 5408 4972 5410 4992
rect 5354 4936 5410 4972
rect 5354 3576 5410 3632
rect 846 2388 848 2408
rect 848 2388 900 2408
rect 900 2388 902 2408
rect 846 2352 902 2388
rect 4802 2252 4804 2272
rect 4804 2252 4856 2272
rect 4856 2252 4858 2272
rect 4802 2216 4858 2252
rect 2616 2202 2672 2204
rect 2696 2202 2752 2204
rect 2776 2202 2832 2204
rect 2856 2202 2912 2204
rect 2616 2150 2662 2202
rect 2662 2150 2672 2202
rect 2696 2150 2726 2202
rect 2726 2150 2738 2202
rect 2738 2150 2752 2202
rect 2776 2150 2790 2202
rect 2790 2150 2802 2202
rect 2802 2150 2832 2202
rect 2856 2150 2866 2202
rect 2866 2150 2912 2202
rect 2616 2148 2672 2150
rect 2696 2148 2752 2150
rect 2776 2148 2832 2150
rect 2856 2148 2912 2150
rect 1674 856 1730 912
rect 5446 856 5502 912
<< metal3 >>
rect 0 10434 800 10464
rect 1393 10434 1459 10437
rect 0 10432 1459 10434
rect 0 10376 1398 10432
rect 1454 10376 1459 10432
rect 0 10374 1459 10376
rect 0 10344 800 10374
rect 1393 10371 1459 10374
rect 4981 10434 5047 10437
rect 6100 10434 6900 10464
rect 4981 10432 6900 10434
rect 4981 10376 4986 10432
rect 5042 10376 6900 10432
rect 4981 10374 6900 10376
rect 4981 10371 5047 10374
rect 6100 10344 6900 10374
rect 1946 9280 2262 9281
rect 1946 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2262 9280
rect 1946 9215 2262 9216
rect 0 9074 800 9104
rect 5349 9074 5415 9077
rect 6100 9074 6900 9104
rect 0 8984 858 9074
rect 5349 9072 6900 9074
rect 5349 9016 5354 9072
rect 5410 9016 6900 9072
rect 5349 9014 6900 9016
rect 5349 9011 5415 9014
rect 6100 8984 6900 9014
rect 798 8941 858 8984
rect 798 8936 907 8941
rect 798 8880 846 8936
rect 902 8880 907 8936
rect 798 8878 907 8880
rect 841 8875 907 8878
rect 2606 8736 2922 8737
rect 2606 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2922 8736
rect 2606 8671 2922 8672
rect 4061 8396 4127 8397
rect 4061 8392 4108 8396
rect 4172 8394 4178 8396
rect 4061 8336 4066 8392
rect 4061 8332 4108 8336
rect 4172 8334 4218 8394
rect 4172 8332 4178 8334
rect 4061 8331 4127 8332
rect 1946 8192 2262 8193
rect 1946 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2262 8192
rect 1946 8127 2262 8128
rect 0 7714 800 7744
rect 933 7714 999 7717
rect 0 7712 999 7714
rect 0 7656 938 7712
rect 994 7656 999 7712
rect 0 7654 999 7656
rect 0 7624 800 7654
rect 933 7651 999 7654
rect 5349 7714 5415 7717
rect 6100 7714 6900 7744
rect 5349 7712 6900 7714
rect 5349 7656 5354 7712
rect 5410 7656 6900 7712
rect 5349 7654 6900 7656
rect 5349 7651 5415 7654
rect 2606 7648 2922 7649
rect 2606 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2922 7648
rect 6100 7624 6900 7654
rect 2606 7583 2922 7584
rect 1946 7104 2262 7105
rect 1946 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2262 7104
rect 1946 7039 2262 7040
rect 2606 6560 2922 6561
rect 2606 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2922 6560
rect 2606 6495 2922 6496
rect 841 6490 907 6493
rect 798 6488 907 6490
rect 798 6432 846 6488
rect 902 6432 907 6488
rect 798 6427 907 6432
rect 798 6384 858 6427
rect 0 6294 858 6384
rect 5349 6354 5415 6357
rect 6100 6354 6900 6384
rect 5349 6352 6900 6354
rect 5349 6296 5354 6352
rect 5410 6296 6900 6352
rect 5349 6294 6900 6296
rect 0 6264 800 6294
rect 5349 6291 5415 6294
rect 6100 6264 6900 6294
rect 1946 6016 2262 6017
rect 1946 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2262 6016
rect 1946 5951 2262 5952
rect 2606 5472 2922 5473
rect 2606 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2922 5472
rect 2606 5407 2922 5408
rect 841 5130 907 5133
rect 798 5128 907 5130
rect 798 5072 846 5128
rect 902 5072 907 5128
rect 798 5067 907 5072
rect 798 5024 858 5067
rect 0 4934 858 5024
rect 5349 4994 5415 4997
rect 6100 4994 6900 5024
rect 5349 4992 6900 4994
rect 5349 4936 5354 4992
rect 5410 4936 6900 4992
rect 5349 4934 6900 4936
rect 0 4904 800 4934
rect 5349 4931 5415 4934
rect 1946 4928 2262 4929
rect 1946 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2262 4928
rect 6100 4904 6900 4934
rect 1946 4863 2262 4864
rect 2606 4384 2922 4385
rect 2606 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2922 4384
rect 2606 4319 2922 4320
rect 4102 3980 4108 4044
rect 4172 4042 4178 4044
rect 4245 4042 4311 4045
rect 4172 4040 4311 4042
rect 4172 3984 4250 4040
rect 4306 3984 4311 4040
rect 4172 3982 4311 3984
rect 4172 3980 4178 3982
rect 4245 3979 4311 3982
rect 1946 3840 2262 3841
rect 1946 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2262 3840
rect 1946 3775 2262 3776
rect 841 3770 907 3773
rect 798 3768 907 3770
rect 798 3712 846 3768
rect 902 3712 907 3768
rect 798 3707 907 3712
rect 798 3664 858 3707
rect 0 3574 858 3664
rect 5349 3634 5415 3637
rect 6100 3634 6900 3664
rect 5349 3632 6900 3634
rect 5349 3576 5354 3632
rect 5410 3576 6900 3632
rect 5349 3574 6900 3576
rect 0 3544 800 3574
rect 5349 3571 5415 3574
rect 6100 3544 6900 3574
rect 2606 3296 2922 3297
rect 2606 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2922 3296
rect 2606 3231 2922 3232
rect 1946 2752 2262 2753
rect 1946 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2262 2752
rect 1946 2687 2262 2688
rect 841 2410 907 2413
rect 798 2408 907 2410
rect 798 2352 846 2408
rect 902 2352 907 2408
rect 798 2347 907 2352
rect 798 2304 858 2347
rect 0 2214 858 2304
rect 4797 2274 4863 2277
rect 6100 2274 6900 2304
rect 4797 2272 6900 2274
rect 4797 2216 4802 2272
rect 4858 2216 6900 2272
rect 4797 2214 6900 2216
rect 0 2184 800 2214
rect 4797 2211 4863 2214
rect 2606 2208 2922 2209
rect 2606 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2922 2208
rect 6100 2184 6900 2214
rect 2606 2143 2922 2144
rect 0 914 800 944
rect 1669 914 1735 917
rect 0 912 1735 914
rect 0 856 1674 912
rect 1730 856 1735 912
rect 0 854 1735 856
rect 0 824 800 854
rect 1669 851 1735 854
rect 5441 914 5507 917
rect 6100 914 6900 944
rect 5441 912 6900 914
rect 5441 856 5446 912
rect 5502 856 6900 912
rect 5441 854 6900 856
rect 5441 851 5507 854
rect 6100 824 6900 854
<< via3 >>
rect 1952 9276 2016 9280
rect 1952 9220 1956 9276
rect 1956 9220 2012 9276
rect 2012 9220 2016 9276
rect 1952 9216 2016 9220
rect 2032 9276 2096 9280
rect 2032 9220 2036 9276
rect 2036 9220 2092 9276
rect 2092 9220 2096 9276
rect 2032 9216 2096 9220
rect 2112 9276 2176 9280
rect 2112 9220 2116 9276
rect 2116 9220 2172 9276
rect 2172 9220 2176 9276
rect 2112 9216 2176 9220
rect 2192 9276 2256 9280
rect 2192 9220 2196 9276
rect 2196 9220 2252 9276
rect 2252 9220 2256 9276
rect 2192 9216 2256 9220
rect 2612 8732 2676 8736
rect 2612 8676 2616 8732
rect 2616 8676 2672 8732
rect 2672 8676 2676 8732
rect 2612 8672 2676 8676
rect 2692 8732 2756 8736
rect 2692 8676 2696 8732
rect 2696 8676 2752 8732
rect 2752 8676 2756 8732
rect 2692 8672 2756 8676
rect 2772 8732 2836 8736
rect 2772 8676 2776 8732
rect 2776 8676 2832 8732
rect 2832 8676 2836 8732
rect 2772 8672 2836 8676
rect 2852 8732 2916 8736
rect 2852 8676 2856 8732
rect 2856 8676 2912 8732
rect 2912 8676 2916 8732
rect 2852 8672 2916 8676
rect 4108 8392 4172 8396
rect 4108 8336 4122 8392
rect 4122 8336 4172 8392
rect 4108 8332 4172 8336
rect 1952 8188 2016 8192
rect 1952 8132 1956 8188
rect 1956 8132 2012 8188
rect 2012 8132 2016 8188
rect 1952 8128 2016 8132
rect 2032 8188 2096 8192
rect 2032 8132 2036 8188
rect 2036 8132 2092 8188
rect 2092 8132 2096 8188
rect 2032 8128 2096 8132
rect 2112 8188 2176 8192
rect 2112 8132 2116 8188
rect 2116 8132 2172 8188
rect 2172 8132 2176 8188
rect 2112 8128 2176 8132
rect 2192 8188 2256 8192
rect 2192 8132 2196 8188
rect 2196 8132 2252 8188
rect 2252 8132 2256 8188
rect 2192 8128 2256 8132
rect 2612 7644 2676 7648
rect 2612 7588 2616 7644
rect 2616 7588 2672 7644
rect 2672 7588 2676 7644
rect 2612 7584 2676 7588
rect 2692 7644 2756 7648
rect 2692 7588 2696 7644
rect 2696 7588 2752 7644
rect 2752 7588 2756 7644
rect 2692 7584 2756 7588
rect 2772 7644 2836 7648
rect 2772 7588 2776 7644
rect 2776 7588 2832 7644
rect 2832 7588 2836 7644
rect 2772 7584 2836 7588
rect 2852 7644 2916 7648
rect 2852 7588 2856 7644
rect 2856 7588 2912 7644
rect 2912 7588 2916 7644
rect 2852 7584 2916 7588
rect 1952 7100 2016 7104
rect 1952 7044 1956 7100
rect 1956 7044 2012 7100
rect 2012 7044 2016 7100
rect 1952 7040 2016 7044
rect 2032 7100 2096 7104
rect 2032 7044 2036 7100
rect 2036 7044 2092 7100
rect 2092 7044 2096 7100
rect 2032 7040 2096 7044
rect 2112 7100 2176 7104
rect 2112 7044 2116 7100
rect 2116 7044 2172 7100
rect 2172 7044 2176 7100
rect 2112 7040 2176 7044
rect 2192 7100 2256 7104
rect 2192 7044 2196 7100
rect 2196 7044 2252 7100
rect 2252 7044 2256 7100
rect 2192 7040 2256 7044
rect 2612 6556 2676 6560
rect 2612 6500 2616 6556
rect 2616 6500 2672 6556
rect 2672 6500 2676 6556
rect 2612 6496 2676 6500
rect 2692 6556 2756 6560
rect 2692 6500 2696 6556
rect 2696 6500 2752 6556
rect 2752 6500 2756 6556
rect 2692 6496 2756 6500
rect 2772 6556 2836 6560
rect 2772 6500 2776 6556
rect 2776 6500 2832 6556
rect 2832 6500 2836 6556
rect 2772 6496 2836 6500
rect 2852 6556 2916 6560
rect 2852 6500 2856 6556
rect 2856 6500 2912 6556
rect 2912 6500 2916 6556
rect 2852 6496 2916 6500
rect 1952 6012 2016 6016
rect 1952 5956 1956 6012
rect 1956 5956 2012 6012
rect 2012 5956 2016 6012
rect 1952 5952 2016 5956
rect 2032 6012 2096 6016
rect 2032 5956 2036 6012
rect 2036 5956 2092 6012
rect 2092 5956 2096 6012
rect 2032 5952 2096 5956
rect 2112 6012 2176 6016
rect 2112 5956 2116 6012
rect 2116 5956 2172 6012
rect 2172 5956 2176 6012
rect 2112 5952 2176 5956
rect 2192 6012 2256 6016
rect 2192 5956 2196 6012
rect 2196 5956 2252 6012
rect 2252 5956 2256 6012
rect 2192 5952 2256 5956
rect 2612 5468 2676 5472
rect 2612 5412 2616 5468
rect 2616 5412 2672 5468
rect 2672 5412 2676 5468
rect 2612 5408 2676 5412
rect 2692 5468 2756 5472
rect 2692 5412 2696 5468
rect 2696 5412 2752 5468
rect 2752 5412 2756 5468
rect 2692 5408 2756 5412
rect 2772 5468 2836 5472
rect 2772 5412 2776 5468
rect 2776 5412 2832 5468
rect 2832 5412 2836 5468
rect 2772 5408 2836 5412
rect 2852 5468 2916 5472
rect 2852 5412 2856 5468
rect 2856 5412 2912 5468
rect 2912 5412 2916 5468
rect 2852 5408 2916 5412
rect 1952 4924 2016 4928
rect 1952 4868 1956 4924
rect 1956 4868 2012 4924
rect 2012 4868 2016 4924
rect 1952 4864 2016 4868
rect 2032 4924 2096 4928
rect 2032 4868 2036 4924
rect 2036 4868 2092 4924
rect 2092 4868 2096 4924
rect 2032 4864 2096 4868
rect 2112 4924 2176 4928
rect 2112 4868 2116 4924
rect 2116 4868 2172 4924
rect 2172 4868 2176 4924
rect 2112 4864 2176 4868
rect 2192 4924 2256 4928
rect 2192 4868 2196 4924
rect 2196 4868 2252 4924
rect 2252 4868 2256 4924
rect 2192 4864 2256 4868
rect 2612 4380 2676 4384
rect 2612 4324 2616 4380
rect 2616 4324 2672 4380
rect 2672 4324 2676 4380
rect 2612 4320 2676 4324
rect 2692 4380 2756 4384
rect 2692 4324 2696 4380
rect 2696 4324 2752 4380
rect 2752 4324 2756 4380
rect 2692 4320 2756 4324
rect 2772 4380 2836 4384
rect 2772 4324 2776 4380
rect 2776 4324 2832 4380
rect 2832 4324 2836 4380
rect 2772 4320 2836 4324
rect 2852 4380 2916 4384
rect 2852 4324 2856 4380
rect 2856 4324 2912 4380
rect 2912 4324 2916 4380
rect 2852 4320 2916 4324
rect 4108 3980 4172 4044
rect 1952 3836 2016 3840
rect 1952 3780 1956 3836
rect 1956 3780 2012 3836
rect 2012 3780 2016 3836
rect 1952 3776 2016 3780
rect 2032 3836 2096 3840
rect 2032 3780 2036 3836
rect 2036 3780 2092 3836
rect 2092 3780 2096 3836
rect 2032 3776 2096 3780
rect 2112 3836 2176 3840
rect 2112 3780 2116 3836
rect 2116 3780 2172 3836
rect 2172 3780 2176 3836
rect 2112 3776 2176 3780
rect 2192 3836 2256 3840
rect 2192 3780 2196 3836
rect 2196 3780 2252 3836
rect 2252 3780 2256 3836
rect 2192 3776 2256 3780
rect 2612 3292 2676 3296
rect 2612 3236 2616 3292
rect 2616 3236 2672 3292
rect 2672 3236 2676 3292
rect 2612 3232 2676 3236
rect 2692 3292 2756 3296
rect 2692 3236 2696 3292
rect 2696 3236 2752 3292
rect 2752 3236 2756 3292
rect 2692 3232 2756 3236
rect 2772 3292 2836 3296
rect 2772 3236 2776 3292
rect 2776 3236 2832 3292
rect 2832 3236 2836 3292
rect 2772 3232 2836 3236
rect 2852 3292 2916 3296
rect 2852 3236 2856 3292
rect 2856 3236 2912 3292
rect 2912 3236 2916 3292
rect 2852 3232 2916 3236
rect 1952 2748 2016 2752
rect 1952 2692 1956 2748
rect 1956 2692 2012 2748
rect 2012 2692 2016 2748
rect 1952 2688 2016 2692
rect 2032 2748 2096 2752
rect 2032 2692 2036 2748
rect 2036 2692 2092 2748
rect 2092 2692 2096 2748
rect 2032 2688 2096 2692
rect 2112 2748 2176 2752
rect 2112 2692 2116 2748
rect 2116 2692 2172 2748
rect 2172 2692 2176 2748
rect 2112 2688 2176 2692
rect 2192 2748 2256 2752
rect 2192 2692 2196 2748
rect 2196 2692 2252 2748
rect 2252 2692 2256 2748
rect 2192 2688 2256 2692
rect 2612 2204 2676 2208
rect 2612 2148 2616 2204
rect 2616 2148 2672 2204
rect 2672 2148 2676 2204
rect 2612 2144 2676 2148
rect 2692 2204 2756 2208
rect 2692 2148 2696 2204
rect 2696 2148 2752 2204
rect 2752 2148 2756 2204
rect 2692 2144 2756 2148
rect 2772 2204 2836 2208
rect 2772 2148 2776 2204
rect 2776 2148 2832 2204
rect 2832 2148 2836 2204
rect 2772 2144 2836 2148
rect 2852 2204 2916 2208
rect 2852 2148 2856 2204
rect 2856 2148 2912 2204
rect 2912 2148 2916 2204
rect 2852 2144 2916 2148
<< metal4 >>
rect 1944 9280 2264 9296
rect 1944 9216 1952 9280
rect 2016 9216 2032 9280
rect 2096 9216 2112 9280
rect 2176 9216 2192 9280
rect 2256 9216 2264 9280
rect 1944 8192 2264 9216
rect 1944 8128 1952 8192
rect 2016 8128 2032 8192
rect 2096 8128 2112 8192
rect 2176 8128 2192 8192
rect 2256 8128 2264 8192
rect 1944 7104 2264 8128
rect 1944 7040 1952 7104
rect 2016 7040 2032 7104
rect 2096 7040 2112 7104
rect 2176 7040 2192 7104
rect 2256 7040 2264 7104
rect 1944 6016 2264 7040
rect 1944 5952 1952 6016
rect 2016 5952 2032 6016
rect 2096 5952 2112 6016
rect 2176 5952 2192 6016
rect 2256 5952 2264 6016
rect 1944 4928 2264 5952
rect 1944 4864 1952 4928
rect 2016 4864 2032 4928
rect 2096 4864 2112 4928
rect 2176 4864 2192 4928
rect 2256 4864 2264 4928
rect 1944 3840 2264 4864
rect 1944 3776 1952 3840
rect 2016 3776 2032 3840
rect 2096 3776 2112 3840
rect 2176 3776 2192 3840
rect 2256 3776 2264 3840
rect 1944 2752 2264 3776
rect 1944 2688 1952 2752
rect 2016 2688 2032 2752
rect 2096 2688 2112 2752
rect 2176 2688 2192 2752
rect 2256 2688 2264 2752
rect 1944 2128 2264 2688
rect 2604 8736 2924 9296
rect 2604 8672 2612 8736
rect 2676 8672 2692 8736
rect 2756 8672 2772 8736
rect 2836 8672 2852 8736
rect 2916 8672 2924 8736
rect 2604 7648 2924 8672
rect 4107 8396 4173 8397
rect 4107 8332 4108 8396
rect 4172 8332 4173 8396
rect 4107 8331 4173 8332
rect 2604 7584 2612 7648
rect 2676 7584 2692 7648
rect 2756 7584 2772 7648
rect 2836 7584 2852 7648
rect 2916 7584 2924 7648
rect 2604 6560 2924 7584
rect 2604 6496 2612 6560
rect 2676 6496 2692 6560
rect 2756 6496 2772 6560
rect 2836 6496 2852 6560
rect 2916 6496 2924 6560
rect 2604 5472 2924 6496
rect 2604 5408 2612 5472
rect 2676 5408 2692 5472
rect 2756 5408 2772 5472
rect 2836 5408 2852 5472
rect 2916 5408 2924 5472
rect 2604 4384 2924 5408
rect 2604 4320 2612 4384
rect 2676 4320 2692 4384
rect 2756 4320 2772 4384
rect 2836 4320 2852 4384
rect 2916 4320 2924 4384
rect 2604 3296 2924 4320
rect 4110 4045 4170 8331
rect 4107 4044 4173 4045
rect 4107 3980 4108 4044
rect 4172 3980 4173 4044
rect 4107 3979 4173 3980
rect 2604 3232 2612 3296
rect 2676 3232 2692 3296
rect 2756 3232 2772 3296
rect 2836 3232 2852 3296
rect 2916 3232 2924 3296
rect 2604 2208 2924 3232
rect 2604 2144 2612 2208
rect 2676 2144 2692 2208
rect 2756 2144 2772 2208
rect 2836 2144 2852 2208
rect 2916 2144 2924 2208
rect 2604 2128 2924 2144
use sky130_fd_sc_hd__nor2_1  _10_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _11_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2300 0 1 5440
box -38 -48 682 592
use sky130_fd_sc_hd__o31a_1  _12_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4876 0 -1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__or4_2  _13_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2668 0 -1 8704
box -38 -48 682 592
use sky130_fd_sc_hd__and2b_1  _14_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4784 0 1 6528
box -38 -48 590 592
use sky130_fd_sc_hd__clkbuf_1  _15_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform -1 0 5152 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__nor2_1  _16_
timestamp 1704896540
transform 1 0 5060 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__and2_1  _17_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 -1 8704
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _18_
timestamp 1704896540
transform 1 0 4232 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__xnor2_1  _19_
timestamp 1704896540
transform 1 0 3772 0 1 2176
box -38 -48 682 592
use sky130_fd_sc_hd__or4_1  _20_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2760 0 -1 5440
box -38 -48 590 592
use sky130_fd_sc_hd__o31ai_1  _21_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 2760 0 1 8704
box -38 -48 590 592
use sky130_fd_sc_hd__and2_1  _22_
timestamp 1704896540
transform 1 0 3864 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__clkbuf_1  _23_
timestamp 1704896540
transform 1 0 4692 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__xor2_1  _24_ $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4508 0 1 3264
box -38 -48 682 592
use sky130_fd_sc_hd__and2_1  _25_
timestamp 1704896540
transform -1 0 3588 0 -1 7616
box -38 -48 498 592
use sky130_fd_sc_hd__nor2_1  _26_
timestamp 1704896540
transform -1 0 1840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  _27_
timestamp 1704896540
transform -1 0 3588 0 -1 8704
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_0_9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1932 0 1 2176
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_0_21 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3036 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_0_27 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3588 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_0_36 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4416 0 1 2176
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_3
timestamp 1704896540
transform 1 0 1380 0 -1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_1_15
timestamp 1704896540
transform 1 0 2484 0 -1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_1_27
timestamp 1704896540
transform 1 0 3588 0 -1 3264
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_1_33
timestamp 1704896540
transform 1 0 4140 0 -1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_1_37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4508 0 -1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_3
timestamp 1704896540
transform 1 0 1380 0 1 3264
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_2_15
timestamp 1704896540
transform 1 0 2484 0 1 3264
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_2_27
timestamp 1704896540
transform 1 0 3588 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_2_29 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3772 0 1 3264
box -38 -48 774 592
use sky130_fd_sc_hd__decap_4  FILLER_0_2_44
timestamp 1704896540
transform 1 0 5152 0 1 3264
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_6
timestamp 1704896540
transform 1 0 1656 0 -1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_3_18
timestamp 1704896540
transform 1 0 2760 0 -1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_3_30
timestamp 1704896540
transform 1 0 3864 0 -1 4352
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_3_38
timestamp 1704896540
transform 1 0 4600 0 -1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_3_42
timestamp 1704896540
transform 1 0 4968 0 -1 4352
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_3
timestamp 1704896540
transform 1 0 1380 0 1 4352
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_15
timestamp 1704896540
transform 1 0 2484 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_27
timestamp 1704896540
transform 1 0 3588 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_4_29
timestamp 1704896540
transform 1 0 3772 0 1 4352
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_4_41
timestamp 1704896540
transform 1 0 4876 0 1 4352
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_4_47
timestamp 1704896540
transform 1 0 5428 0 1 4352
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_6
timestamp 1704896540
transform 1 0 1656 0 -1 5440
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_5_24
timestamp 1704896540
transform 1 0 3312 0 -1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_5_36
timestamp 1704896540
transform 1 0 4416 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_5_40
timestamp 1704896540
transform 1 0 4784 0 -1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_3
timestamp 1704896540
transform 1 0 1380 0 1 5440
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_6_11
timestamp 1704896540
transform 1 0 2116 0 1 5440
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_6_20
timestamp 1704896540
transform 1 0 2944 0 1 5440
box -38 -48 774 592
use sky130_ef_sc_hd__decap_12  FILLER_0_6_32
timestamp 1704896540
transform 1 0 4048 0 1 5440
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_6_44
timestamp 1704896540
transform 1 0 5152 0 1 5440
box -38 -48 406 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_3
timestamp 1704896540
transform 1 0 1380 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_15
timestamp 1704896540
transform 1 0 2484 0 -1 6528
box -38 -48 1142 592
use sky130_ef_sc_hd__decap_12  FILLER_0_7_27
timestamp 1704896540
transform 1 0 3588 0 -1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_7_39
timestamp 1704896540
transform 1 0 4692 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_7_43
timestamp 1704896540
transform 1 0 5060 0 -1 6528
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_8_6
timestamp 1704896540
transform 1 0 1656 0 1 6528
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_18
timestamp 1704896540
transform 1 0 2760 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_26
timestamp 1704896540
transform 1 0 3496 0 1 6528
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_8_29
timestamp 1704896540
transform 1 0 3772 0 1 6528
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_8_37 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4508 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__fill_2  FILLER_0_8_46
timestamp 1704896540
transform 1 0 5336 0 1 6528
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_3
timestamp 1704896540
transform 1 0 1380 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_6  FILLER_0_9_15
timestamp 1704896540
transform 1 0 2484 0 -1 7616
box -38 -48 590 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_21
timestamp 1704896540
transform 1 0 3036 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__decap_3  FILLER_0_9_27
timestamp 1704896540
transform 1 0 3588 0 -1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_9_35
timestamp 1704896540
transform 1 0 4324 0 -1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_1  FILLER_0_9_47
timestamp 1704896540
transform 1 0 5428 0 -1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__fill_2  FILLER_0_10_3
timestamp 1704896540
transform 1 0 1380 0 1 7616
box -38 -48 222 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_11
timestamp 1704896540
transform 1 0 2116 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_4  FILLER_0_10_23
timestamp 1704896540
transform 1 0 3220 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__fill_1  FILLER_0_10_27
timestamp 1704896540
transform 1 0 3588 0 1 7616
box -38 -48 130 592
use sky130_ef_sc_hd__decap_12  FILLER_0_10_29
timestamp 1704896540
transform 1 0 3772 0 1 7616
box -38 -48 1142 592
use sky130_fd_sc_hd__decap_3  FILLER_0_10_41
timestamp 1704896540
transform 1 0 4876 0 1 7616
box -38 -48 314 592
use sky130_ef_sc_hd__decap_12  FILLER_0_11_3
timestamp 1704896540
transform 1 0 1380 0 -1 8704
box -38 -48 1142 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_15
timestamp 1704896540
transform 1 0 2484 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_1  FILLER_0_11_27
timestamp 1704896540
transform 1 0 3588 0 -1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_8  FILLER_0_11_33
timestamp 1704896540
transform 1 0 4140 0 -1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_41
timestamp 1704896540
transform 1 0 4876 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__fill_2  FILLER_0_11_46
timestamp 1704896540
transform 1 0 5336 0 -1 8704
box -38 -48 222 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_9
timestamp 1704896540
transform 1 0 1932 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__fill_1  FILLER_0_12_17
timestamp 1704896540
transform 1 0 2668 0 1 8704
box -38 -48 130 592
use sky130_fd_sc_hd__decap_4  FILLER_0_12_24
timestamp 1704896540
transform 1 0 3312 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__decap_8  FILLER_0_12_29
timestamp 1704896540
transform 1 0 3772 0 1 8704
box -38 -48 774 592
use sky130_fd_sc_hd__decap_3  FILLER_0_12_37
timestamp 1704896540
transform 1 0 4508 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input1 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 1380 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input2
timestamp 1704896540
transform 1 0 1656 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input3
timestamp 1704896540
transform 1 0 1840 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input4
timestamp 1704896540
transform 1 0 1380 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input5
timestamp 1704896540
transform 1 0 1380 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input6
timestamp 1704896540
transform 1 0 1380 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__buf_1  input7
timestamp 1704896540
transform 1 0 1380 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__clkbuf_1  input8
timestamp 1704896540
transform -1 0 1932 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__buf_2  output9 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4784 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output10
timestamp 1704896540
transform 1 0 5152 0 1 8704
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output11
timestamp 1704896540
transform 1 0 5152 0 1 7616
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output12
timestamp 1704896540
transform 1 0 5152 0 -1 6528
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output13
timestamp 1704896540
transform 1 0 5152 0 -1 5440
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output14
timestamp 1704896540
transform 1 0 5152 0 -1 4352
box -38 -48 406 592
use sky130_fd_sc_hd__buf_2  output15
timestamp 1704896540
transform 1 0 4600 0 1 2176
box -38 -48 406 592
use sky130_fd_sc_hd__clkbuf_4  output16 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 4968 0 1 2176
box -38 -48 590 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Left_13
timestamp 1704896540
transform 1 0 1104 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_0_Right_0
timestamp 1704896540
transform -1 0 5796 0 1 2176
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Left_14
timestamp 1704896540
transform 1 0 1104 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_1_Right_1
timestamp 1704896540
transform -1 0 5796 0 -1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Left_15
timestamp 1704896540
transform 1 0 1104 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_2_Right_2
timestamp 1704896540
transform -1 0 5796 0 1 3264
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Left_16
timestamp 1704896540
transform 1 0 1104 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_3_Right_3
timestamp 1704896540
transform -1 0 5796 0 -1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Left_17
timestamp 1704896540
transform 1 0 1104 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_4_Right_4
timestamp 1704896540
transform -1 0 5796 0 1 4352
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Left_18
timestamp 1704896540
transform 1 0 1104 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_5_Right_5
timestamp 1704896540
transform -1 0 5796 0 -1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Left_19
timestamp 1704896540
transform 1 0 1104 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_6_Right_6
timestamp 1704896540
transform -1 0 5796 0 1 5440
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Left_20
timestamp 1704896540
transform 1 0 1104 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_7_Right_7
timestamp 1704896540
transform -1 0 5796 0 -1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Left_21
timestamp 1704896540
transform 1 0 1104 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_8_Right_8
timestamp 1704896540
transform -1 0 5796 0 1 6528
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Left_22
timestamp 1704896540
transform 1 0 1104 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_9_Right_9
timestamp 1704896540
transform -1 0 5796 0 -1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Left_23
timestamp 1704896540
transform 1 0 1104 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_10_Right_10
timestamp 1704896540
transform -1 0 5796 0 1 7616
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Left_24
timestamp 1704896540
transform 1 0 1104 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_11_Right_11
timestamp 1704896540
transform -1 0 5796 0 -1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Left_25
timestamp 1704896540
transform 1 0 1104 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__decap_3  PHY_EDGE_ROW_12_Right_12
timestamp 1704896540
transform -1 0 5796 0 1 8704
box -38 -48 314 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_0_26 $PDKPATH/libs.ref/sky130_fd_sc_hd/mag
timestamp 1704896540
transform 1 0 3680 0 1 2176
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_2_27
timestamp 1704896540
transform 1 0 3680 0 1 3264
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_4_28
timestamp 1704896540
transform 1 0 3680 0 1 4352
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_6_29
timestamp 1704896540
transform 1 0 3680 0 1 5440
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_8_30
timestamp 1704896540
transform 1 0 3680 0 1 6528
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_10_31
timestamp 1704896540
transform 1 0 3680 0 1 7616
box -38 -48 130 592
use sky130_fd_sc_hd__tapvpwrvgnd_1  TAP_TAPCELL_ROW_12_32
timestamp 1704896540
transform 1 0 3680 0 1 8704
box -38 -48 130 592
<< labels >>
flabel metal4 s 2604 2128 2924 9296 0 FreeSans 1920 90 0 0 VGND
port 0 nsew ground bidirectional
flabel metal4 s 1944 2128 2264 9296 0 FreeSans 1920 90 0 0 VPWR
port 1 nsew power bidirectional
flabel metal3 s 0 10344 800 10464 0 FreeSans 480 0 0 0 in[0]
port 2 nsew signal input
flabel metal3 s 0 8984 800 9104 0 FreeSans 480 0 0 0 in[1]
port 3 nsew signal input
flabel metal3 s 0 7624 800 7744 0 FreeSans 480 0 0 0 in[2]
port 4 nsew signal input
flabel metal3 s 0 6264 800 6384 0 FreeSans 480 0 0 0 in[3]
port 5 nsew signal input
flabel metal3 s 0 4904 800 5024 0 FreeSans 480 0 0 0 in[4]
port 6 nsew signal input
flabel metal3 s 0 3544 800 3664 0 FreeSans 480 0 0 0 in[5]
port 7 nsew signal input
flabel metal3 s 0 2184 800 2304 0 FreeSans 480 0 0 0 in[6]
port 8 nsew signal input
flabel metal3 s 0 824 800 944 0 FreeSans 480 0 0 0 in[7]
port 9 nsew signal input
flabel metal3 s 6100 10344 6900 10464 0 FreeSans 480 0 0 0 out[0]
port 10 nsew signal output
flabel metal3 s 6100 8984 6900 9104 0 FreeSans 480 0 0 0 out[1]
port 11 nsew signal output
flabel metal3 s 6100 7624 6900 7744 0 FreeSans 480 0 0 0 out[2]
port 12 nsew signal output
flabel metal3 s 6100 6264 6900 6384 0 FreeSans 480 0 0 0 out[3]
port 13 nsew signal output
flabel metal3 s 6100 4904 6900 5024 0 FreeSans 480 0 0 0 out[4]
port 14 nsew signal output
flabel metal3 s 6100 3544 6900 3664 0 FreeSans 480 0 0 0 out[5]
port 15 nsew signal output
flabel metal3 s 6100 2184 6900 2304 0 FreeSans 480 0 0 0 out[6]
port 16 nsew signal output
flabel metal3 s 6100 824 6900 944 0 FreeSans 480 0 0 0 out[7]
port 17 nsew signal output
rlabel metal1 3450 8704 3450 8704 0 VGND
rlabel metal1 3450 9248 3450 9248 0 VPWR
rlabel metal1 2024 5746 2024 5746 0 _00_
rlabel metal1 4876 3162 4876 3162 0 _01_
rlabel metal1 3588 5066 3588 5066 0 _02_
rlabel metal2 4922 5916 4922 5916 0 _03_
rlabel metal1 4278 2482 4278 2482 0 _04_
rlabel metal3 4209 4012 4209 4012 0 _05_
rlabel metal2 3266 4284 3266 4284 0 _06_
rlabel metal1 4048 7378 4048 7378 0 _07_
rlabel metal1 4600 4114 4600 4114 0 _08_
rlabel metal1 2484 7514 2484 7514 0 _09_
rlabel metal3 1050 10404 1050 10404 0 in[0]
rlabel metal3 751 9044 751 9044 0 in[1]
rlabel metal3 820 7684 820 7684 0 in[2]
rlabel metal3 751 6324 751 6324 0 in[3]
rlabel metal3 751 4964 751 4964 0 in[4]
rlabel metal3 751 3604 751 3604 0 in[5]
rlabel metal3 751 2244 751 2244 0 in[6]
rlabel metal3 1188 884 1188 884 0 in[7]
rlabel metal2 3818 4284 3818 4284 0 net1
rlabel metal1 3496 7990 3496 7990 0 net10
rlabel metal1 3542 5814 3542 5814 0 net11
rlabel metal1 5152 5338 5152 5338 0 net12
rlabel metal1 4692 3094 4692 3094 0 net13
rlabel metal1 4784 2550 4784 2550 0 net14
rlabel metal2 4646 3162 4646 3162 0 net15
rlabel metal2 5106 2992 5106 2992 0 net16
rlabel metal2 4002 4318 4002 4318 0 net2
rlabel metal1 2530 5644 2530 5644 0 net3
rlabel metal1 2392 6630 2392 6630 0 net4
rlabel metal1 3220 5202 3220 5202 0 net5
rlabel metal2 3082 3706 3082 3706 0 net6
rlabel metal2 2990 3842 2990 3842 0 net7
rlabel metal1 3312 2618 3312 2618 0 net8
rlabel metal2 3542 8772 3542 8772 0 net9
rlabel metal2 5014 9775 5014 9775 0 out[0]
rlabel via2 5382 9061 5382 9061 0 out[1]
rlabel via2 5382 7701 5382 7701 0 out[2]
rlabel metal2 5382 6375 5382 6375 0 out[3]
rlabel via2 5382 4981 5382 4981 0 out[4]
rlabel metal2 5382 3757 5382 3757 0 out[5]
rlabel via2 4830 2261 4830 2261 0 out[6]
rlabel metal2 5474 1615 5474 1615 0 out[7]
<< properties >>
string FIXED_BBOX 0 0 6900 11424
<< end >>
